magic
tech scmos
timestamp 1731999991
<< nwell >>
rect 187 53 257 77
rect 267 53 303 77
rect 267 41 331 53
rect 307 27 331 41
rect 187 -34 268 -10
rect 284 -51 328 -41
rect 284 -77 357 -51
rect 187 -129 257 -105
rect 187 -218 275 -194
rect 284 -242 336 -225
rect 284 -261 371 -242
rect 339 -268 371 -261
rect 187 -316 268 -292
rect 187 -409 257 -385
<< ntransistor >>
rect 198 20 200 32
rect 210 20 212 32
rect 241 20 243 26
rect 280 11 282 17
rect 288 11 290 17
rect 318 11 320 17
rect 198 -74 200 -62
rect 210 -74 212 -62
rect 222 -74 224 -62
rect 252 -71 254 -65
rect 344 -93 346 -87
rect 297 -114 299 -108
rect 305 -114 307 -108
rect 313 -114 315 -108
rect 198 -162 200 -150
rect 210 -162 212 -150
rect 241 -162 243 -156
rect 198 -265 200 -253
rect 210 -265 212 -253
rect 222 -265 224 -253
rect 234 -265 236 -253
rect 259 -262 261 -256
rect 358 -284 360 -278
rect 297 -306 299 -300
rect 305 -306 307 -300
rect 313 -306 315 -300
rect 321 -306 323 -300
rect 198 -356 200 -344
rect 210 -356 212 -344
rect 222 -356 224 -344
rect 252 -353 254 -347
rect 198 -442 200 -430
rect 210 -442 212 -430
rect 241 -442 243 -436
<< ptransistor >>
rect 198 59 200 71
rect 210 59 212 71
rect 241 59 243 71
rect 280 47 282 71
rect 288 47 290 71
rect 318 33 320 45
rect 198 -28 200 -16
rect 210 -28 212 -16
rect 222 -28 224 -16
rect 252 -28 254 -16
rect 297 -71 299 -47
rect 305 -71 307 -47
rect 313 -71 315 -47
rect 344 -71 346 -59
rect 198 -123 200 -111
rect 210 -123 212 -111
rect 241 -123 243 -111
rect 198 -212 200 -200
rect 210 -212 212 -200
rect 222 -212 224 -200
rect 234 -212 236 -200
rect 259 -212 261 -200
rect 297 -255 299 -231
rect 305 -255 307 -231
rect 313 -255 315 -231
rect 321 -255 323 -231
rect 198 -310 200 -298
rect 210 -310 212 -298
rect 222 -310 224 -298
rect 252 -310 254 -298
rect 358 -262 360 -250
rect 198 -403 200 -391
rect 210 -403 212 -391
rect 241 -403 243 -391
<< ndiffusion >>
rect 194 20 198 32
rect 200 20 210 32
rect 212 20 215 32
rect 237 20 241 26
rect 243 20 247 26
rect 277 11 280 17
rect 282 11 283 17
rect 287 11 288 17
rect 290 11 293 17
rect 317 11 318 17
rect 320 11 321 17
rect 194 -74 198 -62
rect 200 -74 210 -62
rect 212 -74 222 -62
rect 224 -74 225 -62
rect 248 -71 252 -65
rect 254 -71 258 -65
rect 343 -93 344 -87
rect 346 -93 347 -87
rect 294 -114 297 -108
rect 299 -114 300 -108
rect 304 -114 305 -108
rect 307 -114 308 -108
rect 312 -114 313 -108
rect 315 -114 318 -108
rect 194 -162 198 -150
rect 200 -162 210 -150
rect 212 -162 215 -150
rect 237 -162 241 -156
rect 243 -162 247 -156
rect 194 -265 198 -253
rect 200 -265 210 -253
rect 212 -265 222 -253
rect 224 -265 234 -253
rect 236 -265 237 -253
rect 255 -262 259 -256
rect 261 -262 265 -256
rect 357 -284 358 -278
rect 360 -284 361 -278
rect 294 -306 297 -300
rect 299 -306 300 -300
rect 304 -306 305 -300
rect 307 -306 308 -300
rect 312 -306 313 -300
rect 315 -306 316 -300
rect 320 -306 321 -300
rect 323 -306 326 -300
rect 194 -356 198 -344
rect 200 -356 210 -344
rect 212 -356 222 -344
rect 224 -356 225 -344
rect 248 -353 252 -347
rect 254 -353 258 -347
rect 194 -442 198 -430
rect 200 -442 210 -430
rect 212 -442 215 -430
rect 237 -442 241 -436
rect 243 -442 247 -436
<< pdiffusion >>
rect 197 59 198 71
rect 200 59 203 71
rect 207 59 210 71
rect 212 59 213 71
rect 237 59 241 71
rect 243 59 247 71
rect 277 47 280 71
rect 282 47 288 71
rect 290 47 293 71
rect 317 33 318 45
rect 320 33 321 45
rect 197 -28 198 -16
rect 200 -28 203 -16
rect 207 -28 210 -16
rect 212 -28 215 -16
rect 219 -28 222 -16
rect 224 -28 225 -16
rect 248 -28 252 -16
rect 254 -28 258 -16
rect 294 -71 297 -47
rect 299 -71 305 -47
rect 307 -71 313 -47
rect 315 -71 318 -47
rect 343 -71 344 -59
rect 346 -71 347 -59
rect 197 -123 198 -111
rect 200 -123 203 -111
rect 207 -123 210 -111
rect 212 -123 213 -111
rect 237 -123 241 -111
rect 243 -123 247 -111
rect 197 -212 198 -200
rect 200 -212 203 -200
rect 207 -212 210 -200
rect 212 -212 215 -200
rect 219 -212 222 -200
rect 224 -212 227 -200
rect 231 -212 234 -200
rect 236 -212 237 -200
rect 255 -212 259 -200
rect 261 -212 265 -200
rect 294 -255 297 -231
rect 299 -255 305 -231
rect 307 -255 313 -231
rect 315 -255 321 -231
rect 323 -255 326 -231
rect 197 -310 198 -298
rect 200 -310 203 -298
rect 207 -310 210 -298
rect 212 -310 215 -298
rect 219 -310 222 -298
rect 224 -310 225 -298
rect 248 -310 252 -298
rect 254 -310 258 -298
rect 357 -262 358 -250
rect 360 -262 361 -250
rect 197 -403 198 -391
rect 200 -403 203 -391
rect 207 -403 210 -391
rect 212 -403 213 -391
rect 237 -403 241 -391
rect 243 -403 247 -391
<< ndcontact >>
rect 190 20 194 32
rect 215 20 219 32
rect 233 20 237 26
rect 247 20 251 26
rect 273 11 277 17
rect 283 11 287 17
rect 293 11 297 17
rect 313 11 317 17
rect 321 11 325 17
rect 190 -74 194 -62
rect 225 -74 229 -62
rect 244 -71 248 -65
rect 258 -71 262 -65
rect 339 -93 343 -87
rect 347 -93 351 -87
rect 290 -114 294 -108
rect 300 -114 304 -108
rect 308 -114 312 -108
rect 318 -114 322 -108
rect 190 -162 194 -150
rect 215 -162 219 -150
rect 233 -162 237 -156
rect 247 -162 251 -156
rect 190 -265 194 -253
rect 237 -265 241 -253
rect 251 -262 255 -256
rect 265 -262 269 -256
rect 353 -284 357 -278
rect 361 -284 365 -278
rect 290 -306 294 -300
rect 300 -306 304 -300
rect 308 -306 312 -300
rect 316 -306 320 -300
rect 326 -306 330 -300
rect 190 -356 194 -344
rect 225 -356 229 -344
rect 244 -353 248 -347
rect 258 -353 262 -347
rect 190 -442 194 -430
rect 215 -442 219 -430
rect 233 -442 237 -436
rect 247 -442 251 -436
<< pdcontact >>
rect 193 59 197 71
rect 203 59 207 71
rect 213 59 217 71
rect 233 59 237 71
rect 247 59 251 71
rect 273 47 277 71
rect 293 47 297 71
rect 313 33 317 45
rect 321 33 325 45
rect 193 -28 197 -16
rect 203 -28 207 -16
rect 215 -28 219 -16
rect 225 -28 229 -16
rect 244 -28 248 -16
rect 258 -28 262 -16
rect 290 -71 294 -47
rect 318 -71 322 -47
rect 339 -71 343 -59
rect 347 -71 351 -59
rect 193 -123 197 -111
rect 203 -123 207 -111
rect 213 -123 217 -111
rect 233 -123 237 -111
rect 247 -123 251 -111
rect 193 -212 197 -200
rect 203 -212 207 -200
rect 215 -212 219 -200
rect 227 -212 231 -200
rect 237 -212 241 -200
rect 251 -212 255 -200
rect 265 -212 269 -200
rect 290 -255 294 -231
rect 326 -255 330 -231
rect 193 -310 197 -298
rect 203 -310 207 -298
rect 215 -310 219 -298
rect 225 -310 229 -298
rect 244 -310 248 -298
rect 258 -310 262 -298
rect 353 -262 357 -250
rect 361 -262 365 -250
rect 193 -403 197 -391
rect 203 -403 207 -391
rect 213 -403 217 -391
rect 233 -403 237 -391
rect 247 -403 251 -391
<< polysilicon >>
rect 198 71 200 74
rect 210 71 212 74
rect 241 71 243 74
rect 280 71 282 74
rect 288 71 290 74
rect 198 32 200 59
rect 210 32 212 59
rect 241 26 243 59
rect 280 38 282 47
rect 198 17 200 20
rect 210 17 212 20
rect 241 17 243 20
rect 280 17 282 34
rect 288 31 290 47
rect 318 45 320 48
rect 288 17 290 27
rect 318 17 320 33
rect 280 8 282 11
rect 288 8 290 11
rect 318 7 320 11
rect 198 -16 200 -13
rect 210 -16 212 -13
rect 222 -16 224 -13
rect 252 -16 254 -13
rect 198 -62 200 -28
rect 210 -62 212 -28
rect 222 -62 224 -28
rect 252 -65 254 -28
rect 297 -47 299 -44
rect 305 -47 307 -44
rect 313 -47 315 -44
rect 344 -59 346 -56
rect 252 -74 254 -71
rect 198 -77 200 -74
rect 210 -77 212 -74
rect 222 -77 224 -74
rect 297 -80 299 -71
rect 297 -108 299 -84
rect 305 -87 307 -71
rect 305 -108 307 -91
rect 313 -94 315 -71
rect 344 -87 346 -71
rect 344 -97 346 -93
rect 313 -108 315 -98
rect 198 -111 200 -108
rect 210 -111 212 -108
rect 241 -111 243 -108
rect 297 -117 299 -114
rect 305 -117 307 -114
rect 313 -117 315 -114
rect 198 -150 200 -123
rect 210 -150 212 -123
rect 241 -156 243 -123
rect 198 -165 200 -162
rect 210 -165 212 -162
rect 241 -165 243 -162
rect 198 -200 200 -197
rect 210 -200 212 -197
rect 222 -200 224 -197
rect 234 -200 236 -197
rect 259 -200 261 -197
rect 198 -253 200 -212
rect 210 -253 212 -212
rect 222 -253 224 -212
rect 234 -253 236 -212
rect 259 -256 261 -212
rect 297 -231 299 -228
rect 305 -231 307 -228
rect 313 -231 315 -228
rect 321 -231 323 -228
rect 358 -250 360 -247
rect 259 -265 261 -262
rect 297 -264 299 -255
rect 198 -268 200 -265
rect 210 -268 212 -265
rect 222 -268 224 -265
rect 234 -268 236 -265
rect 198 -298 200 -295
rect 210 -298 212 -295
rect 222 -298 224 -295
rect 252 -298 254 -295
rect 297 -300 299 -268
rect 305 -271 307 -255
rect 305 -300 307 -275
rect 313 -278 315 -255
rect 313 -300 315 -282
rect 321 -285 323 -255
rect 358 -278 360 -262
rect 358 -288 360 -284
rect 321 -300 323 -289
rect 297 -309 299 -306
rect 305 -309 307 -306
rect 313 -309 315 -306
rect 321 -309 323 -306
rect 198 -344 200 -310
rect 210 -344 212 -310
rect 222 -344 224 -310
rect 252 -347 254 -310
rect 252 -356 254 -353
rect 198 -359 200 -356
rect 210 -359 212 -356
rect 222 -359 224 -356
rect 198 -391 200 -388
rect 210 -391 212 -388
rect 241 -391 243 -388
rect 198 -430 200 -403
rect 210 -430 212 -403
rect 241 -436 243 -403
rect 198 -445 200 -442
rect 210 -445 212 -442
rect 241 -445 243 -442
<< polycontact >>
rect 194 42 198 46
rect 206 35 210 39
rect 237 46 241 50
rect 278 34 282 38
rect 286 27 290 31
rect 314 20 318 24
rect 194 -45 198 -41
rect 206 -52 210 -48
rect 218 -59 222 -55
rect 248 -41 252 -37
rect 295 -84 299 -80
rect 303 -91 307 -87
rect 340 -84 344 -80
rect 311 -98 315 -94
rect 194 -140 198 -136
rect 206 -147 210 -143
rect 237 -136 241 -132
rect 194 -229 198 -225
rect 206 -236 210 -232
rect 218 -243 222 -239
rect 230 -250 234 -246
rect 255 -225 259 -221
rect 295 -268 299 -264
rect 303 -275 307 -271
rect 311 -282 315 -278
rect 354 -275 358 -271
rect 319 -289 323 -285
rect 194 -327 198 -323
rect 206 -334 210 -330
rect 218 -341 222 -337
rect 248 -323 252 -319
rect 194 -420 198 -416
rect 206 -427 210 -423
rect 237 -416 241 -412
<< metal1 >>
rect 187 75 237 79
rect 267 75 306 79
rect 193 71 197 75
rect 213 71 217 75
rect 233 71 237 75
rect 273 71 277 75
rect 203 50 207 59
rect 247 50 251 59
rect 203 46 237 50
rect 247 46 264 50
rect 302 53 306 75
rect 302 49 317 53
rect 149 42 194 46
rect 149 -55 153 42
rect 156 35 206 39
rect 156 -45 160 35
rect 215 32 219 46
rect 247 26 251 46
rect 260 38 264 46
rect 260 34 278 38
rect 260 27 286 31
rect 190 15 194 20
rect 233 15 237 20
rect 187 11 237 15
rect 260 8 264 27
rect 293 24 297 47
rect 313 45 317 49
rect 321 24 325 33
rect 283 20 314 24
rect 321 20 329 24
rect 283 17 287 20
rect 321 17 325 20
rect 164 4 264 8
rect 273 7 277 11
rect 293 7 297 11
rect 313 7 317 11
rect 164 -36 168 4
rect 267 3 317 7
rect 187 -12 248 -8
rect 193 -16 197 -12
rect 215 -16 219 -12
rect 244 -16 248 -12
rect 203 -37 207 -28
rect 225 -37 229 -28
rect 258 -37 262 -28
rect 203 -41 248 -37
rect 258 -41 281 -37
rect 161 -48 174 -45
rect 161 -49 206 -48
rect 170 -52 206 -49
rect 149 -59 218 -55
rect 149 -246 153 -59
rect 225 -62 229 -41
rect 156 -239 160 -69
rect 165 -143 169 -68
rect 258 -65 262 -41
rect 190 -79 194 -74
rect 244 -79 248 -71
rect 187 -83 248 -79
rect 277 -80 281 -41
rect 284 -43 329 -39
rect 290 -47 294 -43
rect 325 -51 329 -43
rect 325 -55 343 -51
rect 339 -59 343 -55
rect 318 -80 322 -71
rect 347 -80 351 -71
rect 277 -84 295 -80
rect 318 -84 340 -80
rect 347 -84 355 -80
rect 260 -91 303 -87
rect 187 -107 237 -103
rect 193 -111 197 -107
rect 213 -111 217 -107
rect 233 -111 237 -107
rect 203 -132 207 -123
rect 247 -132 251 -123
rect 260 -132 264 -91
rect 203 -136 237 -132
rect 247 -136 264 -132
rect 276 -98 311 -94
rect 165 -147 206 -143
rect 165 -226 169 -147
rect 215 -150 219 -136
rect 247 -156 251 -136
rect 190 -167 194 -162
rect 233 -167 237 -162
rect 187 -171 237 -167
rect 276 -174 280 -98
rect 318 -101 322 -84
rect 347 -87 351 -84
rect 339 -97 343 -93
rect 300 -105 322 -101
rect 300 -108 304 -105
rect 318 -108 322 -105
rect 325 -101 343 -97
rect 290 -118 294 -114
rect 308 -118 312 -114
rect 325 -118 329 -101
rect 284 -122 329 -118
rect 173 -178 280 -174
rect 173 -209 177 -178
rect 187 -196 255 -192
rect 193 -200 197 -196
rect 215 -200 219 -196
rect 237 -200 241 -196
rect 251 -200 255 -196
rect 203 -221 207 -212
rect 227 -221 231 -212
rect 265 -221 269 -212
rect 203 -225 255 -221
rect 265 -225 281 -221
rect 174 -229 194 -225
rect 156 -243 218 -239
rect 149 -250 230 -246
rect 237 -253 241 -225
rect 152 -423 156 -259
rect 164 -337 168 -259
rect 173 -323 177 -259
rect 265 -256 269 -225
rect 190 -270 194 -265
rect 251 -270 255 -262
rect 277 -264 281 -225
rect 284 -227 338 -223
rect 290 -231 294 -227
rect 334 -242 338 -227
rect 334 -246 357 -242
rect 277 -268 295 -264
rect 187 -274 255 -270
rect 326 -271 330 -255
rect 353 -250 357 -246
rect 361 -271 365 -262
rect 270 -275 303 -271
rect 326 -275 354 -271
rect 361 -275 369 -271
rect 187 -294 248 -290
rect 193 -298 197 -294
rect 215 -298 219 -294
rect 244 -298 248 -294
rect 203 -319 207 -310
rect 225 -319 229 -310
rect 258 -319 262 -310
rect 270 -319 274 -275
rect 309 -282 311 -278
rect 203 -323 248 -319
rect 258 -323 274 -319
rect 277 -289 319 -285
rect 173 -327 194 -323
rect 173 -328 177 -327
rect 164 -341 218 -337
rect 225 -344 229 -323
rect 172 -416 176 -350
rect 258 -347 262 -323
rect 190 -361 194 -356
rect 244 -361 248 -353
rect 187 -365 248 -361
rect 187 -387 237 -383
rect 193 -391 197 -387
rect 213 -391 217 -387
rect 233 -391 237 -387
rect 203 -412 207 -403
rect 247 -412 251 -403
rect 277 -412 281 -289
rect 326 -293 330 -275
rect 361 -278 365 -275
rect 353 -288 357 -284
rect 300 -297 330 -293
rect 339 -292 357 -288
rect 300 -300 304 -297
rect 316 -300 320 -297
rect 290 -310 294 -306
rect 308 -310 312 -306
rect 326 -310 330 -306
rect 339 -310 343 -292
rect 284 -314 343 -310
rect 203 -416 237 -412
rect 247 -416 281 -412
rect 172 -420 194 -416
rect 152 -427 206 -423
rect 215 -430 219 -416
rect 247 -436 251 -416
rect 190 -447 194 -442
rect 233 -447 237 -442
rect 187 -451 237 -447
<< m2contact >>
rect 164 -41 169 -36
rect 156 -50 161 -45
rect 156 -69 161 -64
rect 165 -68 170 -63
rect 173 -214 178 -209
rect 164 -231 169 -226
rect 173 -234 178 -229
rect 152 -259 157 -254
rect 163 -259 168 -254
rect 173 -259 178 -254
rect 172 -333 177 -328
rect 172 -350 177 -345
<< metal2 >>
rect 156 -64 160 -50
rect 165 -63 169 -41
rect 185 -45 194 -41
rect 185 -136 189 -45
rect 185 -140 194 -136
rect 173 -218 177 -214
rect 152 -222 177 -218
rect 152 -254 156 -222
rect 164 -254 168 -231
rect 174 -254 178 -234
rect 185 -232 189 -140
rect 185 -236 206 -232
rect 185 -330 189 -236
rect 172 -345 176 -333
rect 185 -334 206 -330
<< labels >>
rlabel metal1 301 -225 301 -225 5 VDD
rlabel pdcontact 292 -243 292 -243 1 vdd
rlabel metal1 302 -312 302 -312 1 GND
rlabel ndcontact 310 -303 310 -303 1 gnd
rlabel ndcontact 292 -303 292 -303 1 gnd
rlabel ndcontact 328 -303 328 -303 1 gnd
rlabel ndcontact 355 -281 355 -281 1 gnd
rlabel pdcontact 355 -256 355 -256 1 vdd
rlabel metal1 205 -292 205 -292 5 VDD
rlabel metal1 192 -363 192 -363 2 GND
rlabel ndcontact 192 -350 192 -350 3 gnd
rlabel ndcontact 246 -350 246 -350 1 gnd
rlabel pdcontact 246 -304 246 -304 1 vdd
rlabel pdcontact 217 -304 217 -304 1 vdd
rlabel pdcontact 195 -304 195 -304 1 vdd
rlabel metal1 205 77 205 77 5 VDD
rlabel metal1 192 13 192 13 2 GND
rlabel metal1 285 5 285 5 1 GND
rlabel metal1 284 77 284 77 5 VDD
rlabel metal1 205 -10 205 -10 5 VDD
rlabel metal1 192 -81 192 -81 2 GND
rlabel ndcontact 192 -68 192 -68 3 gnd
rlabel ndcontact 246 -68 246 -68 1 gnd
rlabel pdcontact 246 -22 246 -22 1 vdd
rlabel pdcontact 217 -22 217 -22 1 vdd
rlabel pdcontact 195 -22 195 -22 1 vdd
rlabel metal1 205 -105 205 -105 5 VDD
rlabel metal1 192 -169 192 -169 2 GND
rlabel metal1 301 -41 301 -41 5 VDD
rlabel metal1 302 -120 302 -120 1 GND
rlabel ndcontact 341 -90 341 -90 1 gnd
rlabel pdcontact 341 -65 341 -65 1 vdd
rlabel ndcontact 310 -111 310 -111 1 gnd
rlabel ndcontact 292 -111 292 -111 1 gnd
rlabel pdcontact 292 -59 292 -59 1 vdd
rlabel metal1 205 -194 205 -194 5 VDD
rlabel pdcontact 217 -206 217 -206 1 vdd
rlabel pdcontact 195 -206 195 -206 1 vdd
rlabel ndcontact 192 -259 192 -259 3 gnd
rlabel metal1 192 -272 192 -272 2 GND
rlabel pdcontact 253 -206 253 -206 1 vdd
rlabel ndcontact 253 -259 253 -259 1 gnd
rlabel pdcontact 239 -206 239 -206 1 vdd
rlabel metal1 205 -385 205 -385 5 VDD
rlabel metal1 192 -449 192 -449 2 GND
rlabel polycontact 196 44 196 44 1 g0
rlabel polycontact 239 48 239 48 1 p1g0_bar
rlabel polycontact 280 36 280 36 1 p1g0
rlabel polycontact 288 29 288 29 1 g1
rlabel polycontact 316 22 316 22 1 c2_bar
rlabel metal1 327 22 327 22 1 c2
rlabel pdcontact 195 65 195 65 1 vdd
rlabel pdcontact 215 65 215 65 1 vdd
rlabel pdcontact 205 65 205 65 1 p1g0_bar
rlabel ndcontact 217 26 217 26 1 p1g0_bar
rlabel ndcontact 192 26 192 26 3 gnd
rlabel pdcontact 235 65 235 65 1 vdd
rlabel pdcontact 249 65 249 65 1 p1g0
rlabel ndcontact 235 23 235 23 1 gnd
rlabel ndcontact 249 23 249 23 1 p1g0
rlabel pdcontact 275 59 275 59 1 vdd
rlabel ndcontact 275 14 275 14 1 gnd
rlabel ndcontact 295 14 295 14 1 gnd
rlabel ndcontact 285 14 285 14 1 c2_bar
rlabel pdcontact 295 59 295 59 1 c2_bar
rlabel ndcontact 315 14 315 14 1 gnd
rlabel ndcontact 323 14 323 14 1 c2
rlabel pdcontact 323 39 323 39 1 c2
rlabel pdcontact 315 39 315 39 1 vdd
rlabel ndiffusion 205 26 205 26 1 n1
rlabel pdiffusion 285 60 285 60 1 n2
rlabel polycontact 220 -57 220 -57 1 g0
rlabel ndiffusion 205 -68 205 -68 1 n3
rlabel ndiffusion 217 -68 217 -68 1 n4
rlabel polycontact 250 -39 250 -39 1 p2p1g0_bar
rlabel pdcontact 227 -22 227 -22 1 p2p1g0_bar
rlabel pdcontact 205 -22 205 -22 1 p2p1g0_bar
rlabel pdcontact 260 -22 260 -22 1 p2p1g0
rlabel ndcontact 260 -68 260 -68 1 p2p1g0
rlabel ndcontact 227 -68 227 -68 1 p2p1g0_bar
rlabel polycontact 297 -82 297 -82 1 p2p1g0
rlabel pdcontact 215 -117 215 -117 1 vdd
rlabel pdcontact 235 -117 235 -117 1 vdd
rlabel pdcontact 195 -117 195 -117 1 vdd
rlabel polycontact 208 -145 208 -145 1 g1
rlabel polycontact 239 -134 239 -134 1 p2g1_bar
rlabel pdcontact 205 -117 205 -117 1 p2g1_bar
rlabel ndcontact 217 -156 217 -156 1 p2g1_bar
rlabel ndcontact 192 -156 192 -156 3 gnd
rlabel ndcontact 235 -159 235 -159 1 gnd
rlabel pdcontact 249 -117 249 -117 1 p2g1
rlabel ndcontact 249 -159 249 -159 1 p2g1
rlabel polycontact 305 -89 305 -89 1 p2g1
rlabel polycontact 313 -96 313 -96 1 g2
rlabel ndcontact 302 -111 302 -111 1 c3_bar
rlabel ndcontact 320 -111 320 -111 1 c3_bar
rlabel pdcontact 320 -59 320 -59 1 c3_bar
rlabel polycontact 342 -82 342 -82 1 c3_bar
rlabel metal1 353 -82 353 -82 1 c3
rlabel ndcontact 349 -90 349 -90 1 c3
rlabel pdcontact 349 -65 349 -65 1 c3
rlabel polycontact 232 -248 232 -248 1 g0
rlabel ndiffusion 205 -156 205 -156 1 n5
rlabel pdiffusion 302 -59 302 -59 1 n6
rlabel pdiffusion 310 -59 310 -59 1 n7
rlabel ndiffusion 205 -259 205 -259 1 n8
rlabel ndiffusion 217 -259 217 -259 1 n9
rlabel ndiffusion 229 -259 229 -259 1 n10
rlabel ndcontact 239 -259 239 -259 1 p3p2p1g0_bar
rlabel pdcontact 229 -206 229 -206 1 p3p2p1g0_bar
rlabel pdcontact 205 -206 205 -206 1 p3p2p1g0_bar
rlabel polycontact 257 -223 257 -223 1 p3p2p1g0_bar
rlabel ndcontact 267 -259 267 -259 1 p3p2p1g0
rlabel pdcontact 267 -206 267 -206 1 p3p2p1g0
rlabel polycontact 297 -266 297 -266 1 p3p2p1g0
rlabel polycontact 220 -339 220 -339 1 g1
rlabel ndiffusion 205 -350 205 -350 1 n11
rlabel ndiffusion 217 -350 217 -350 1 n12
rlabel ndcontact 227 -350 227 -350 1 p3p2g1_bar
rlabel pdcontact 205 -304 205 -304 1 p3p2g1_bar
rlabel pdcontact 227 -304 227 -304 1 p3p2g1_bar
rlabel polycontact 250 -321 250 -321 1 p3p2g1_bar
rlabel ndcontact 260 -350 260 -350 1 p3p2g1
rlabel pdcontact 260 -304 260 -304 1 p3p2g1
rlabel polycontact 305 -273 305 -273 1 p3p2g1
rlabel polycontact 208 -425 208 -425 1 g2
rlabel ndcontact 192 -436 192 -436 3 gnd
rlabel ndcontact 235 -439 235 -439 1 gnd
rlabel ndcontact 217 -436 217 -436 1 p3g2_bar
rlabel pdcontact 195 -397 195 -397 1 vdd
rlabel pdcontact 205 -397 205 -397 1 p3g2_bar
rlabel pdcontact 215 -397 215 -397 1 vdd
rlabel polycontact 239 -414 239 -414 1 p3g2_bar
rlabel pdcontact 235 -397 235 -397 1 vdd
rlabel pdcontact 249 -397 249 -397 1 p3g2
rlabel ndcontact 249 -439 249 -439 1 p3g2
rlabel ndiffusion 205 -436 205 -436 1 n13
rlabel polycontact 321 -287 321 -287 1 p3g2
rlabel pdiffusion 302 -242 302 -242 1 n14
rlabel pdiffusion 310 -242 310 -242 1 n15
rlabel pdiffusion 318 -242 318 -242 1 n16
rlabel polycontact 313 -280 313 -280 1 g3
rlabel ndcontact 302 -303 302 -303 1 cout_bar
rlabel ndcontact 318 -303 318 -303 1 cout_bar
rlabel pdcontact 328 -243 328 -243 1 cout_bar
rlabel polycontact 356 -273 356 -273 1 cout_bar
rlabel metal1 367 -273 367 -273 7 cout
rlabel ndcontact 363 -281 363 -281 1 cout
rlabel pdcontact 363 -256 363 -256 1 cout
rlabel polycontact 208 37 208 37 1 p1
rlabel polycontact 208 -50 208 -50 1 p1
rlabel polycontact 220 -241 220 -241 1 p1
rlabel polycontact 196 -43 196 -43 1 p2
rlabel polycontact 196 -138 196 -138 1 p2
rlabel polycontact 208 -234 208 -234 1 p2
rlabel polycontact 208 -332 208 -332 1 p2
rlabel polycontact 196 -227 196 -227 1 p3
rlabel polycontact 196 -325 196 -325 1 p3
rlabel polycontact 196 -418 196 -418 1 p3
<< end >>
