magic
tech scmos
timestamp 1732022920
<< nwell >>
rect 794 631 818 655
rect 828 649 898 673
rect 913 614 949 638
rect 1313 616 1337 640
rect 1347 634 1417 658
rect 913 602 977 614
rect 794 571 818 595
rect 828 571 898 595
rect 953 588 977 602
rect 1432 599 1468 623
rect 1074 564 1144 588
rect 1154 564 1190 588
rect 1432 587 1496 599
rect 906 532 977 556
rect 1154 552 1218 564
rect 1313 556 1337 580
rect 1347 556 1417 580
rect 1472 573 1496 587
rect 1194 538 1218 552
rect 794 469 818 493
rect 828 487 898 511
rect 1074 477 1155 501
rect 910 452 946 476
rect 1171 460 1215 470
rect 910 440 974 452
rect 794 409 818 433
rect 828 409 898 433
rect 950 426 974 440
rect 1171 434 1244 460
rect 1313 452 1337 476
rect 1347 470 1417 494
rect 1432 435 1468 459
rect 1432 423 1496 435
rect 903 370 974 394
rect 1074 382 1144 406
rect 1313 392 1337 416
rect 1347 392 1417 416
rect 1472 409 1496 423
rect 794 307 818 331
rect 828 325 898 349
rect 913 290 949 314
rect 1074 293 1162 317
rect 913 278 977 290
rect 794 247 818 271
rect 828 247 898 271
rect 953 264 977 278
rect 1171 269 1223 286
rect 1313 285 1337 309
rect 1347 303 1417 327
rect 1171 250 1258 269
rect 1432 268 1468 292
rect 1432 256 1496 268
rect 1226 243 1258 250
rect 906 208 977 232
rect 1313 225 1337 249
rect 1347 225 1417 249
rect 1472 242 1496 256
rect 1074 195 1155 219
rect 794 145 818 169
rect 828 163 898 187
rect 910 128 946 152
rect 910 116 974 128
rect 794 85 818 109
rect 828 85 898 109
rect 950 102 974 116
rect 1074 102 1144 126
rect 1314 120 1338 144
rect 1348 138 1418 162
rect 1433 103 1469 127
rect 1433 91 1497 103
rect 903 46 974 70
rect 1314 60 1338 84
rect 1348 60 1418 84
rect 1473 77 1497 91
<< ntransistor >>
rect 805 615 807 621
rect 839 616 841 628
rect 851 616 853 628
rect 882 616 884 622
rect 1324 600 1326 606
rect 1358 601 1360 613
rect 1370 601 1372 613
rect 1401 601 1403 607
rect 805 555 807 561
rect 839 538 841 550
rect 851 538 853 550
rect 926 572 928 578
rect 934 572 936 578
rect 964 572 966 578
rect 882 538 884 544
rect 917 499 919 511
rect 929 499 931 511
rect 1085 531 1087 543
rect 1097 531 1099 543
rect 1128 531 1130 537
rect 1324 540 1326 546
rect 1167 522 1169 528
rect 1175 522 1177 528
rect 1205 522 1207 528
rect 1358 523 1360 535
rect 1370 523 1372 535
rect 1445 557 1447 563
rect 1453 557 1455 563
rect 1483 557 1485 563
rect 1401 523 1403 529
rect 960 499 962 505
rect 805 453 807 459
rect 839 454 841 466
rect 851 454 853 466
rect 882 454 884 460
rect 1085 437 1087 449
rect 1097 437 1099 449
rect 1109 437 1111 449
rect 1139 440 1141 446
rect 805 393 807 399
rect 839 376 841 388
rect 851 376 853 388
rect 923 410 925 416
rect 931 410 933 416
rect 961 410 963 416
rect 1324 436 1326 442
rect 1358 437 1360 449
rect 1370 437 1372 449
rect 1401 437 1403 443
rect 1231 418 1233 424
rect 1184 397 1186 403
rect 1192 397 1194 403
rect 1200 397 1202 403
rect 882 376 884 382
rect 914 337 916 349
rect 926 337 928 349
rect 1085 349 1087 361
rect 1097 349 1099 361
rect 1324 376 1326 382
rect 1358 359 1360 371
rect 1370 359 1372 371
rect 1445 393 1447 399
rect 1453 393 1455 399
rect 1483 393 1485 399
rect 1401 359 1403 365
rect 1128 349 1130 355
rect 957 337 959 343
rect 805 291 807 297
rect 839 292 841 304
rect 851 292 853 304
rect 882 292 884 298
rect 805 231 807 237
rect 839 214 841 226
rect 851 214 853 226
rect 926 248 928 254
rect 934 248 936 254
rect 964 248 966 254
rect 1085 246 1087 258
rect 1097 246 1099 258
rect 1109 246 1111 258
rect 1121 246 1123 258
rect 1324 269 1326 275
rect 1358 270 1360 282
rect 1370 270 1372 282
rect 1401 270 1403 276
rect 1146 249 1148 255
rect 882 214 884 220
rect 917 175 919 187
rect 929 175 931 187
rect 1245 227 1247 233
rect 1184 205 1186 211
rect 1192 205 1194 211
rect 1200 205 1202 211
rect 1208 205 1210 211
rect 1324 209 1326 215
rect 960 175 962 181
rect 805 129 807 135
rect 839 130 841 142
rect 851 130 853 142
rect 1085 155 1087 167
rect 1097 155 1099 167
rect 1109 155 1111 167
rect 1358 192 1360 204
rect 1370 192 1372 204
rect 1445 226 1447 232
rect 1453 226 1455 232
rect 1483 226 1485 232
rect 1401 192 1403 198
rect 1139 158 1141 164
rect 882 130 884 136
rect 805 69 807 75
rect 839 52 841 64
rect 851 52 853 64
rect 923 86 925 92
rect 931 86 933 92
rect 961 86 963 92
rect 1085 69 1087 81
rect 1097 69 1099 81
rect 1325 104 1327 110
rect 1359 105 1361 117
rect 1371 105 1373 117
rect 1402 105 1404 111
rect 1128 69 1130 75
rect 882 52 884 58
rect 914 13 916 25
rect 926 13 928 25
rect 1325 44 1327 50
rect 1359 27 1361 39
rect 1371 27 1373 39
rect 1446 61 1448 67
rect 1454 61 1456 67
rect 1484 61 1486 67
rect 1402 27 1404 33
rect 957 13 959 19
<< ptransistor >>
rect 839 655 841 667
rect 851 655 853 667
rect 882 655 884 667
rect 805 637 807 649
rect 1358 640 1360 652
rect 1370 640 1372 652
rect 1401 640 1403 652
rect 926 608 928 632
rect 934 608 936 632
rect 1324 622 1326 634
rect 805 577 807 589
rect 839 577 841 589
rect 851 577 853 589
rect 882 577 884 589
rect 964 594 966 606
rect 1445 593 1447 617
rect 1453 593 1455 617
rect 1085 570 1087 582
rect 1097 570 1099 582
rect 1128 570 1130 582
rect 917 538 919 550
rect 929 538 931 550
rect 960 538 962 550
rect 839 493 841 505
rect 851 493 853 505
rect 882 493 884 505
rect 1167 558 1169 582
rect 1175 558 1177 582
rect 1324 562 1326 574
rect 1358 562 1360 574
rect 1370 562 1372 574
rect 1401 562 1403 574
rect 1483 579 1485 591
rect 1205 544 1207 556
rect 805 475 807 487
rect 1085 483 1087 495
rect 1097 483 1099 495
rect 1109 483 1111 495
rect 1139 483 1141 495
rect 923 446 925 470
rect 931 446 933 470
rect 805 415 807 427
rect 839 415 841 427
rect 851 415 853 427
rect 882 415 884 427
rect 961 432 963 444
rect 1358 476 1360 488
rect 1370 476 1372 488
rect 1401 476 1403 488
rect 1184 440 1186 464
rect 1192 440 1194 464
rect 1200 440 1202 464
rect 1324 458 1326 470
rect 1231 440 1233 452
rect 1445 429 1447 453
rect 1453 429 1455 453
rect 1085 388 1087 400
rect 1097 388 1099 400
rect 1128 388 1130 400
rect 1324 398 1326 410
rect 1358 398 1360 410
rect 1370 398 1372 410
rect 1401 398 1403 410
rect 1483 415 1485 427
rect 914 376 916 388
rect 926 376 928 388
rect 957 376 959 388
rect 839 331 841 343
rect 851 331 853 343
rect 882 331 884 343
rect 805 313 807 325
rect 926 284 928 308
rect 934 284 936 308
rect 1085 299 1087 311
rect 1097 299 1099 311
rect 1109 299 1111 311
rect 1121 299 1123 311
rect 1146 299 1148 311
rect 1358 309 1360 321
rect 1370 309 1372 321
rect 1401 309 1403 321
rect 805 253 807 265
rect 839 253 841 265
rect 851 253 853 265
rect 882 253 884 265
rect 964 270 966 282
rect 1324 291 1326 303
rect 1184 256 1186 280
rect 1192 256 1194 280
rect 1200 256 1202 280
rect 1208 256 1210 280
rect 1445 262 1447 286
rect 1453 262 1455 286
rect 917 214 919 226
rect 929 214 931 226
rect 960 214 962 226
rect 839 169 841 181
rect 851 169 853 181
rect 882 169 884 181
rect 1085 201 1087 213
rect 1097 201 1099 213
rect 1109 201 1111 213
rect 1139 201 1141 213
rect 1245 249 1247 261
rect 1324 231 1326 243
rect 1358 231 1360 243
rect 1370 231 1372 243
rect 1401 231 1403 243
rect 1483 248 1485 260
rect 805 151 807 163
rect 923 122 925 146
rect 931 122 933 146
rect 1359 144 1361 156
rect 1371 144 1373 156
rect 1402 144 1404 156
rect 1325 126 1327 138
rect 805 91 807 103
rect 839 91 841 103
rect 851 91 853 103
rect 882 91 884 103
rect 961 108 963 120
rect 1085 108 1087 120
rect 1097 108 1099 120
rect 1128 108 1130 120
rect 1446 97 1448 121
rect 1454 97 1456 121
rect 1325 66 1327 78
rect 1359 66 1361 78
rect 1371 66 1373 78
rect 1402 66 1404 78
rect 1484 83 1486 95
rect 914 52 916 64
rect 926 52 928 64
rect 957 52 959 64
<< ndiffusion >>
rect 804 615 805 621
rect 807 615 808 621
rect 835 616 839 628
rect 841 616 851 628
rect 853 616 856 628
rect 878 616 882 622
rect 884 616 888 622
rect 1323 600 1324 606
rect 1326 600 1327 606
rect 1354 601 1358 613
rect 1360 601 1370 613
rect 1372 601 1375 613
rect 1397 601 1401 607
rect 1403 601 1407 607
rect 804 555 805 561
rect 807 555 808 561
rect 835 538 839 550
rect 841 538 851 550
rect 853 538 856 550
rect 923 572 926 578
rect 928 572 929 578
rect 933 572 934 578
rect 936 572 939 578
rect 963 572 964 578
rect 966 572 967 578
rect 878 538 882 544
rect 884 538 888 544
rect 913 499 917 511
rect 919 499 929 511
rect 931 499 934 511
rect 1081 531 1085 543
rect 1087 531 1097 543
rect 1099 531 1102 543
rect 1124 531 1128 537
rect 1130 531 1134 537
rect 1323 540 1324 546
rect 1326 540 1327 546
rect 1164 522 1167 528
rect 1169 522 1170 528
rect 1174 522 1175 528
rect 1177 522 1180 528
rect 1204 522 1205 528
rect 1207 522 1208 528
rect 1354 523 1358 535
rect 1360 523 1370 535
rect 1372 523 1375 535
rect 1442 557 1445 563
rect 1447 557 1448 563
rect 1452 557 1453 563
rect 1455 557 1458 563
rect 1482 557 1483 563
rect 1485 557 1486 563
rect 1397 523 1401 529
rect 1403 523 1407 529
rect 956 499 960 505
rect 962 499 966 505
rect 804 453 805 459
rect 807 453 808 459
rect 835 454 839 466
rect 841 454 851 466
rect 853 454 856 466
rect 878 454 882 460
rect 884 454 888 460
rect 1081 437 1085 449
rect 1087 437 1097 449
rect 1099 437 1109 449
rect 1111 437 1112 449
rect 1135 440 1139 446
rect 1141 440 1145 446
rect 804 393 805 399
rect 807 393 808 399
rect 835 376 839 388
rect 841 376 851 388
rect 853 376 856 388
rect 920 410 923 416
rect 925 410 926 416
rect 930 410 931 416
rect 933 410 936 416
rect 960 410 961 416
rect 963 410 964 416
rect 1323 436 1324 442
rect 1326 436 1327 442
rect 1354 437 1358 449
rect 1360 437 1370 449
rect 1372 437 1375 449
rect 1397 437 1401 443
rect 1403 437 1407 443
rect 1230 418 1231 424
rect 1233 418 1234 424
rect 1181 397 1184 403
rect 1186 397 1187 403
rect 1191 397 1192 403
rect 1194 397 1195 403
rect 1199 397 1200 403
rect 1202 397 1205 403
rect 878 376 882 382
rect 884 376 888 382
rect 910 337 914 349
rect 916 337 926 349
rect 928 337 931 349
rect 1081 349 1085 361
rect 1087 349 1097 361
rect 1099 349 1102 361
rect 1323 376 1324 382
rect 1326 376 1327 382
rect 1354 359 1358 371
rect 1360 359 1370 371
rect 1372 359 1375 371
rect 1442 393 1445 399
rect 1447 393 1448 399
rect 1452 393 1453 399
rect 1455 393 1458 399
rect 1482 393 1483 399
rect 1485 393 1486 399
rect 1397 359 1401 365
rect 1403 359 1407 365
rect 1124 349 1128 355
rect 1130 349 1134 355
rect 953 337 957 343
rect 959 337 963 343
rect 804 291 805 297
rect 807 291 808 297
rect 835 292 839 304
rect 841 292 851 304
rect 853 292 856 304
rect 878 292 882 298
rect 884 292 888 298
rect 804 231 805 237
rect 807 231 808 237
rect 835 214 839 226
rect 841 214 851 226
rect 853 214 856 226
rect 923 248 926 254
rect 928 248 929 254
rect 933 248 934 254
rect 936 248 939 254
rect 963 248 964 254
rect 966 248 967 254
rect 1081 246 1085 258
rect 1087 246 1097 258
rect 1099 246 1109 258
rect 1111 246 1121 258
rect 1123 246 1124 258
rect 1323 269 1324 275
rect 1326 269 1327 275
rect 1354 270 1358 282
rect 1360 270 1370 282
rect 1372 270 1375 282
rect 1397 270 1401 276
rect 1403 270 1407 276
rect 1142 249 1146 255
rect 1148 249 1152 255
rect 878 214 882 220
rect 884 214 888 220
rect 913 175 917 187
rect 919 175 929 187
rect 931 175 934 187
rect 1244 227 1245 233
rect 1247 227 1248 233
rect 1181 205 1184 211
rect 1186 205 1187 211
rect 1191 205 1192 211
rect 1194 205 1195 211
rect 1199 205 1200 211
rect 1202 205 1203 211
rect 1207 205 1208 211
rect 1210 205 1213 211
rect 1323 209 1324 215
rect 1326 209 1327 215
rect 956 175 960 181
rect 962 175 966 181
rect 804 129 805 135
rect 807 129 808 135
rect 835 130 839 142
rect 841 130 851 142
rect 853 130 856 142
rect 1081 155 1085 167
rect 1087 155 1097 167
rect 1099 155 1109 167
rect 1111 155 1112 167
rect 1354 192 1358 204
rect 1360 192 1370 204
rect 1372 192 1375 204
rect 1442 226 1445 232
rect 1447 226 1448 232
rect 1452 226 1453 232
rect 1455 226 1458 232
rect 1482 226 1483 232
rect 1485 226 1486 232
rect 1397 192 1401 198
rect 1403 192 1407 198
rect 1135 158 1139 164
rect 1141 158 1145 164
rect 878 130 882 136
rect 884 130 888 136
rect 804 69 805 75
rect 807 69 808 75
rect 835 52 839 64
rect 841 52 851 64
rect 853 52 856 64
rect 920 86 923 92
rect 925 86 926 92
rect 930 86 931 92
rect 933 86 936 92
rect 960 86 961 92
rect 963 86 964 92
rect 1081 69 1085 81
rect 1087 69 1097 81
rect 1099 69 1102 81
rect 1324 104 1325 110
rect 1327 104 1328 110
rect 1355 105 1359 117
rect 1361 105 1371 117
rect 1373 105 1376 117
rect 1398 105 1402 111
rect 1404 105 1408 111
rect 1124 69 1128 75
rect 1130 69 1134 75
rect 878 52 882 58
rect 884 52 888 58
rect 910 13 914 25
rect 916 13 926 25
rect 928 13 931 25
rect 1324 44 1325 50
rect 1327 44 1328 50
rect 1355 27 1359 39
rect 1361 27 1371 39
rect 1373 27 1376 39
rect 1443 61 1446 67
rect 1448 61 1449 67
rect 1453 61 1454 67
rect 1456 61 1459 67
rect 1483 61 1484 67
rect 1486 61 1487 67
rect 1398 27 1402 33
rect 1404 27 1408 33
rect 953 13 957 19
rect 959 13 963 19
<< pdiffusion >>
rect 838 655 839 667
rect 841 655 844 667
rect 848 655 851 667
rect 853 655 854 667
rect 878 655 882 667
rect 884 655 888 667
rect 804 637 805 649
rect 807 637 808 649
rect 1357 640 1358 652
rect 1360 640 1363 652
rect 1367 640 1370 652
rect 1372 640 1373 652
rect 1397 640 1401 652
rect 1403 640 1407 652
rect 923 608 926 632
rect 928 608 934 632
rect 936 608 939 632
rect 1323 622 1324 634
rect 1326 622 1327 634
rect 804 577 805 589
rect 807 577 808 589
rect 838 577 839 589
rect 841 577 844 589
rect 848 577 851 589
rect 853 577 854 589
rect 878 577 882 589
rect 884 577 888 589
rect 963 594 964 606
rect 966 594 967 606
rect 1442 593 1445 617
rect 1447 593 1453 617
rect 1455 593 1458 617
rect 1084 570 1085 582
rect 1087 570 1090 582
rect 1094 570 1097 582
rect 1099 570 1100 582
rect 1124 570 1128 582
rect 1130 570 1134 582
rect 916 538 917 550
rect 919 538 922 550
rect 926 538 929 550
rect 931 538 932 550
rect 956 538 960 550
rect 962 538 966 550
rect 838 493 839 505
rect 841 493 844 505
rect 848 493 851 505
rect 853 493 854 505
rect 878 493 882 505
rect 884 493 888 505
rect 1164 558 1167 582
rect 1169 558 1175 582
rect 1177 558 1180 582
rect 1323 562 1324 574
rect 1326 562 1327 574
rect 1357 562 1358 574
rect 1360 562 1363 574
rect 1367 562 1370 574
rect 1372 562 1373 574
rect 1397 562 1401 574
rect 1403 562 1407 574
rect 1482 579 1483 591
rect 1485 579 1486 591
rect 1204 544 1205 556
rect 1207 544 1208 556
rect 804 475 805 487
rect 807 475 808 487
rect 1084 483 1085 495
rect 1087 483 1090 495
rect 1094 483 1097 495
rect 1099 483 1102 495
rect 1106 483 1109 495
rect 1111 483 1112 495
rect 1135 483 1139 495
rect 1141 483 1145 495
rect 920 446 923 470
rect 925 446 931 470
rect 933 446 936 470
rect 804 415 805 427
rect 807 415 808 427
rect 838 415 839 427
rect 841 415 844 427
rect 848 415 851 427
rect 853 415 854 427
rect 878 415 882 427
rect 884 415 888 427
rect 960 432 961 444
rect 963 432 964 444
rect 1357 476 1358 488
rect 1360 476 1363 488
rect 1367 476 1370 488
rect 1372 476 1373 488
rect 1397 476 1401 488
rect 1403 476 1407 488
rect 1181 440 1184 464
rect 1186 440 1192 464
rect 1194 440 1200 464
rect 1202 440 1205 464
rect 1323 458 1324 470
rect 1326 458 1327 470
rect 1230 440 1231 452
rect 1233 440 1234 452
rect 1442 429 1445 453
rect 1447 429 1453 453
rect 1455 429 1458 453
rect 1084 388 1085 400
rect 1087 388 1090 400
rect 1094 388 1097 400
rect 1099 388 1100 400
rect 1124 388 1128 400
rect 1130 388 1134 400
rect 1323 398 1324 410
rect 1326 398 1327 410
rect 1357 398 1358 410
rect 1360 398 1363 410
rect 1367 398 1370 410
rect 1372 398 1373 410
rect 1397 398 1401 410
rect 1403 398 1407 410
rect 1482 415 1483 427
rect 1485 415 1486 427
rect 913 376 914 388
rect 916 376 919 388
rect 923 376 926 388
rect 928 376 929 388
rect 953 376 957 388
rect 959 376 963 388
rect 838 331 839 343
rect 841 331 844 343
rect 848 331 851 343
rect 853 331 854 343
rect 878 331 882 343
rect 884 331 888 343
rect 804 313 805 325
rect 807 313 808 325
rect 923 284 926 308
rect 928 284 934 308
rect 936 284 939 308
rect 1084 299 1085 311
rect 1087 299 1090 311
rect 1094 299 1097 311
rect 1099 299 1102 311
rect 1106 299 1109 311
rect 1111 299 1114 311
rect 1118 299 1121 311
rect 1123 299 1124 311
rect 1142 299 1146 311
rect 1148 299 1152 311
rect 1357 309 1358 321
rect 1360 309 1363 321
rect 1367 309 1370 321
rect 1372 309 1373 321
rect 1397 309 1401 321
rect 1403 309 1407 321
rect 804 253 805 265
rect 807 253 808 265
rect 838 253 839 265
rect 841 253 844 265
rect 848 253 851 265
rect 853 253 854 265
rect 878 253 882 265
rect 884 253 888 265
rect 963 270 964 282
rect 966 270 967 282
rect 1323 291 1324 303
rect 1326 291 1327 303
rect 1181 256 1184 280
rect 1186 256 1192 280
rect 1194 256 1200 280
rect 1202 256 1208 280
rect 1210 256 1213 280
rect 1442 262 1445 286
rect 1447 262 1453 286
rect 1455 262 1458 286
rect 916 214 917 226
rect 919 214 922 226
rect 926 214 929 226
rect 931 214 932 226
rect 956 214 960 226
rect 962 214 966 226
rect 838 169 839 181
rect 841 169 844 181
rect 848 169 851 181
rect 853 169 854 181
rect 878 169 882 181
rect 884 169 888 181
rect 1084 201 1085 213
rect 1087 201 1090 213
rect 1094 201 1097 213
rect 1099 201 1102 213
rect 1106 201 1109 213
rect 1111 201 1112 213
rect 1135 201 1139 213
rect 1141 201 1145 213
rect 1244 249 1245 261
rect 1247 249 1248 261
rect 1323 231 1324 243
rect 1326 231 1327 243
rect 1357 231 1358 243
rect 1360 231 1363 243
rect 1367 231 1370 243
rect 1372 231 1373 243
rect 1397 231 1401 243
rect 1403 231 1407 243
rect 1482 248 1483 260
rect 1485 248 1486 260
rect 804 151 805 163
rect 807 151 808 163
rect 920 122 923 146
rect 925 122 931 146
rect 933 122 936 146
rect 1358 144 1359 156
rect 1361 144 1364 156
rect 1368 144 1371 156
rect 1373 144 1374 156
rect 1398 144 1402 156
rect 1404 144 1408 156
rect 1324 126 1325 138
rect 1327 126 1328 138
rect 804 91 805 103
rect 807 91 808 103
rect 838 91 839 103
rect 841 91 844 103
rect 848 91 851 103
rect 853 91 854 103
rect 878 91 882 103
rect 884 91 888 103
rect 960 108 961 120
rect 963 108 964 120
rect 1084 108 1085 120
rect 1087 108 1090 120
rect 1094 108 1097 120
rect 1099 108 1100 120
rect 1124 108 1128 120
rect 1130 108 1134 120
rect 1443 97 1446 121
rect 1448 97 1454 121
rect 1456 97 1459 121
rect 1324 66 1325 78
rect 1327 66 1328 78
rect 1358 66 1359 78
rect 1361 66 1364 78
rect 1368 66 1371 78
rect 1373 66 1374 78
rect 1398 66 1402 78
rect 1404 66 1408 78
rect 1483 83 1484 95
rect 1486 83 1487 95
rect 913 52 914 64
rect 916 52 919 64
rect 923 52 926 64
rect 928 52 929 64
rect 953 52 957 64
rect 959 52 963 64
<< ndcontact >>
rect 800 615 804 621
rect 808 615 812 621
rect 831 616 835 628
rect 856 616 860 628
rect 874 616 878 622
rect 888 616 892 622
rect 1319 600 1323 606
rect 1327 600 1331 606
rect 1350 601 1354 613
rect 1375 601 1379 613
rect 1393 601 1397 607
rect 1407 601 1411 607
rect 800 555 804 561
rect 808 555 812 561
rect 831 538 835 550
rect 856 538 860 550
rect 919 572 923 578
rect 929 572 933 578
rect 939 572 943 578
rect 959 572 963 578
rect 967 572 971 578
rect 874 538 878 544
rect 888 538 892 544
rect 909 499 913 511
rect 934 499 938 511
rect 1077 531 1081 543
rect 1102 531 1106 543
rect 1120 531 1124 537
rect 1134 531 1138 537
rect 1319 540 1323 546
rect 1327 540 1331 546
rect 1160 522 1164 528
rect 1170 522 1174 528
rect 1180 522 1184 528
rect 1200 522 1204 528
rect 1208 522 1212 528
rect 1350 523 1354 535
rect 1375 523 1379 535
rect 1438 557 1442 563
rect 1448 557 1452 563
rect 1458 557 1462 563
rect 1478 557 1482 563
rect 1486 557 1490 563
rect 1393 523 1397 529
rect 1407 523 1411 529
rect 952 499 956 505
rect 966 499 970 505
rect 800 453 804 459
rect 808 453 812 459
rect 831 454 835 466
rect 856 454 860 466
rect 874 454 878 460
rect 888 454 892 460
rect 1077 437 1081 449
rect 1112 437 1116 449
rect 1131 440 1135 446
rect 1145 440 1149 446
rect 800 393 804 399
rect 808 393 812 399
rect 831 376 835 388
rect 856 376 860 388
rect 916 410 920 416
rect 926 410 930 416
rect 936 410 940 416
rect 956 410 960 416
rect 964 410 968 416
rect 1319 436 1323 442
rect 1327 436 1331 442
rect 1350 437 1354 449
rect 1375 437 1379 449
rect 1393 437 1397 443
rect 1407 437 1411 443
rect 1226 418 1230 424
rect 1234 418 1238 424
rect 1177 397 1181 403
rect 1187 397 1191 403
rect 1195 397 1199 403
rect 1205 397 1209 403
rect 874 376 878 382
rect 888 376 892 382
rect 906 337 910 349
rect 931 337 935 349
rect 1077 349 1081 361
rect 1102 349 1106 361
rect 1319 376 1323 382
rect 1327 376 1331 382
rect 1350 359 1354 371
rect 1375 359 1379 371
rect 1438 393 1442 399
rect 1448 393 1452 399
rect 1458 393 1462 399
rect 1478 393 1482 399
rect 1486 393 1490 399
rect 1393 359 1397 365
rect 1407 359 1411 365
rect 1120 349 1124 355
rect 1134 349 1138 355
rect 949 337 953 343
rect 963 337 967 343
rect 800 291 804 297
rect 808 291 812 297
rect 831 292 835 304
rect 856 292 860 304
rect 874 292 878 298
rect 888 292 892 298
rect 800 231 804 237
rect 808 231 812 237
rect 831 214 835 226
rect 856 214 860 226
rect 919 248 923 254
rect 929 248 933 254
rect 939 248 943 254
rect 959 248 963 254
rect 967 248 971 254
rect 1077 246 1081 258
rect 1124 246 1128 258
rect 1319 269 1323 275
rect 1327 269 1331 275
rect 1350 270 1354 282
rect 1375 270 1379 282
rect 1393 270 1397 276
rect 1407 270 1411 276
rect 1138 249 1142 255
rect 1152 249 1156 255
rect 874 214 878 220
rect 888 214 892 220
rect 909 175 913 187
rect 934 175 938 187
rect 1240 227 1244 233
rect 1248 227 1252 233
rect 1177 205 1181 211
rect 1187 205 1191 211
rect 1195 205 1199 211
rect 1203 205 1207 211
rect 1213 205 1217 211
rect 1319 209 1323 215
rect 1327 209 1331 215
rect 952 175 956 181
rect 966 175 970 181
rect 800 129 804 135
rect 808 129 812 135
rect 831 130 835 142
rect 856 130 860 142
rect 1077 155 1081 167
rect 1112 155 1116 167
rect 1350 192 1354 204
rect 1375 192 1379 204
rect 1438 226 1442 232
rect 1448 226 1452 232
rect 1458 226 1462 232
rect 1478 226 1482 232
rect 1486 226 1490 232
rect 1393 192 1397 198
rect 1407 192 1411 198
rect 1131 158 1135 164
rect 1145 158 1149 164
rect 874 130 878 136
rect 888 130 892 136
rect 800 69 804 75
rect 808 69 812 75
rect 831 52 835 64
rect 856 52 860 64
rect 916 86 920 92
rect 926 86 930 92
rect 936 86 940 92
rect 956 86 960 92
rect 964 86 968 92
rect 1077 69 1081 81
rect 1102 69 1106 81
rect 1320 104 1324 110
rect 1328 104 1332 110
rect 1351 105 1355 117
rect 1376 105 1380 117
rect 1394 105 1398 111
rect 1408 105 1412 111
rect 1120 69 1124 75
rect 1134 69 1138 75
rect 874 52 878 58
rect 888 52 892 58
rect 906 13 910 25
rect 931 13 935 25
rect 1320 44 1324 50
rect 1328 44 1332 50
rect 1351 27 1355 39
rect 1376 27 1380 39
rect 1439 61 1443 67
rect 1449 61 1453 67
rect 1459 61 1463 67
rect 1479 61 1483 67
rect 1487 61 1491 67
rect 1394 27 1398 33
rect 1408 27 1412 33
rect 949 13 953 19
rect 963 13 967 19
<< pdcontact >>
rect 834 655 838 667
rect 844 655 848 667
rect 854 655 858 667
rect 874 655 878 667
rect 888 655 892 667
rect 800 637 804 649
rect 808 637 812 649
rect 1353 640 1357 652
rect 1363 640 1367 652
rect 1373 640 1377 652
rect 1393 640 1397 652
rect 1407 640 1411 652
rect 919 608 923 632
rect 939 608 943 632
rect 1319 622 1323 634
rect 1327 622 1331 634
rect 800 577 804 589
rect 808 577 812 589
rect 834 577 838 589
rect 844 577 848 589
rect 854 577 858 589
rect 874 577 878 589
rect 888 577 892 589
rect 959 594 963 606
rect 967 594 971 606
rect 1438 593 1442 617
rect 1458 593 1462 617
rect 1080 570 1084 582
rect 1090 570 1094 582
rect 1100 570 1104 582
rect 1120 570 1124 582
rect 1134 570 1138 582
rect 912 538 916 550
rect 922 538 926 550
rect 932 538 936 550
rect 952 538 956 550
rect 966 538 970 550
rect 834 493 838 505
rect 844 493 848 505
rect 854 493 858 505
rect 874 493 878 505
rect 888 493 892 505
rect 1160 558 1164 582
rect 1180 558 1184 582
rect 1319 562 1323 574
rect 1327 562 1331 574
rect 1353 562 1357 574
rect 1363 562 1367 574
rect 1373 562 1377 574
rect 1393 562 1397 574
rect 1407 562 1411 574
rect 1478 579 1482 591
rect 1486 579 1490 591
rect 1200 544 1204 556
rect 1208 544 1212 556
rect 800 475 804 487
rect 808 475 812 487
rect 1080 483 1084 495
rect 1090 483 1094 495
rect 1102 483 1106 495
rect 1112 483 1116 495
rect 1131 483 1135 495
rect 1145 483 1149 495
rect 916 446 920 470
rect 936 446 940 470
rect 800 415 804 427
rect 808 415 812 427
rect 834 415 838 427
rect 844 415 848 427
rect 854 415 858 427
rect 874 415 878 427
rect 888 415 892 427
rect 956 432 960 444
rect 964 432 968 444
rect 1353 476 1357 488
rect 1363 476 1367 488
rect 1373 476 1377 488
rect 1393 476 1397 488
rect 1407 476 1411 488
rect 1177 440 1181 464
rect 1205 440 1209 464
rect 1319 458 1323 470
rect 1327 458 1331 470
rect 1226 440 1230 452
rect 1234 440 1238 452
rect 1438 429 1442 453
rect 1458 429 1462 453
rect 1080 388 1084 400
rect 1090 388 1094 400
rect 1100 388 1104 400
rect 1120 388 1124 400
rect 1134 388 1138 400
rect 1319 398 1323 410
rect 1327 398 1331 410
rect 1353 398 1357 410
rect 1363 398 1367 410
rect 1373 398 1377 410
rect 1393 398 1397 410
rect 1407 398 1411 410
rect 1478 415 1482 427
rect 1486 415 1490 427
rect 909 376 913 388
rect 919 376 923 388
rect 929 376 933 388
rect 949 376 953 388
rect 963 376 967 388
rect 834 331 838 343
rect 844 331 848 343
rect 854 331 858 343
rect 874 331 878 343
rect 888 331 892 343
rect 800 313 804 325
rect 808 313 812 325
rect 919 284 923 308
rect 939 284 943 308
rect 1080 299 1084 311
rect 1090 299 1094 311
rect 1102 299 1106 311
rect 1114 299 1118 311
rect 1124 299 1128 311
rect 1138 299 1142 311
rect 1152 299 1156 311
rect 1353 309 1357 321
rect 1363 309 1367 321
rect 1373 309 1377 321
rect 1393 309 1397 321
rect 1407 309 1411 321
rect 800 253 804 265
rect 808 253 812 265
rect 834 253 838 265
rect 844 253 848 265
rect 854 253 858 265
rect 874 253 878 265
rect 888 253 892 265
rect 959 270 963 282
rect 967 270 971 282
rect 1319 291 1323 303
rect 1327 291 1331 303
rect 1177 256 1181 280
rect 1213 256 1217 280
rect 1438 262 1442 286
rect 1458 262 1462 286
rect 912 214 916 226
rect 922 214 926 226
rect 932 214 936 226
rect 952 214 956 226
rect 966 214 970 226
rect 834 169 838 181
rect 844 169 848 181
rect 854 169 858 181
rect 874 169 878 181
rect 888 169 892 181
rect 1080 201 1084 213
rect 1090 201 1094 213
rect 1102 201 1106 213
rect 1112 201 1116 213
rect 1131 201 1135 213
rect 1145 201 1149 213
rect 1240 249 1244 261
rect 1248 249 1252 261
rect 1319 231 1323 243
rect 1327 231 1331 243
rect 1353 231 1357 243
rect 1363 231 1367 243
rect 1373 231 1377 243
rect 1393 231 1397 243
rect 1407 231 1411 243
rect 1478 248 1482 260
rect 1486 248 1490 260
rect 800 151 804 163
rect 808 151 812 163
rect 916 122 920 146
rect 936 122 940 146
rect 1354 144 1358 156
rect 1364 144 1368 156
rect 1374 144 1378 156
rect 1394 144 1398 156
rect 1408 144 1412 156
rect 1320 126 1324 138
rect 1328 126 1332 138
rect 800 91 804 103
rect 808 91 812 103
rect 834 91 838 103
rect 844 91 848 103
rect 854 91 858 103
rect 874 91 878 103
rect 888 91 892 103
rect 956 108 960 120
rect 964 108 968 120
rect 1080 108 1084 120
rect 1090 108 1094 120
rect 1100 108 1104 120
rect 1120 108 1124 120
rect 1134 108 1138 120
rect 1439 97 1443 121
rect 1459 97 1463 121
rect 1320 66 1324 78
rect 1328 66 1332 78
rect 1354 66 1358 78
rect 1364 66 1368 78
rect 1374 66 1378 78
rect 1394 66 1398 78
rect 1408 66 1412 78
rect 1479 83 1483 95
rect 1487 83 1491 95
rect 909 52 913 64
rect 919 52 923 64
rect 929 52 933 64
rect 949 52 953 64
rect 963 52 967 64
<< polysilicon >>
rect 839 667 841 670
rect 851 667 853 670
rect 882 667 884 670
rect 805 649 807 652
rect 805 621 807 637
rect 839 628 841 655
rect 851 628 853 655
rect 882 622 884 655
rect 1358 652 1360 655
rect 1370 652 1372 655
rect 1401 652 1403 655
rect 926 632 928 635
rect 934 632 936 635
rect 1324 634 1326 637
rect 805 612 807 615
rect 839 613 841 616
rect 851 613 853 616
rect 882 613 884 616
rect 926 599 928 608
rect 805 589 807 592
rect 839 589 841 592
rect 851 589 853 592
rect 882 589 884 592
rect 926 578 928 595
rect 934 592 936 608
rect 964 606 966 609
rect 1324 606 1326 622
rect 1358 613 1360 640
rect 1370 613 1372 640
rect 1401 607 1403 640
rect 1445 617 1447 620
rect 1453 617 1455 620
rect 1324 597 1326 600
rect 1358 598 1360 601
rect 1370 598 1372 601
rect 1401 598 1403 601
rect 934 578 936 588
rect 964 578 966 594
rect 1085 582 1087 585
rect 1097 582 1099 585
rect 1128 582 1130 585
rect 1167 582 1169 585
rect 1175 582 1177 585
rect 1445 584 1447 593
rect 805 561 807 577
rect 805 552 807 555
rect 839 550 841 577
rect 851 550 853 577
rect 882 544 884 577
rect 926 569 928 572
rect 934 569 936 572
rect 964 568 966 572
rect 917 550 919 553
rect 929 550 931 553
rect 960 550 962 553
rect 1085 543 1087 570
rect 1097 543 1099 570
rect 839 535 841 538
rect 851 535 853 538
rect 882 535 884 538
rect 917 511 919 538
rect 929 511 931 538
rect 839 505 841 508
rect 851 505 853 508
rect 882 505 884 508
rect 960 505 962 538
rect 1128 537 1130 570
rect 1324 574 1326 577
rect 1358 574 1360 577
rect 1370 574 1372 577
rect 1401 574 1403 577
rect 1445 563 1447 580
rect 1453 577 1455 593
rect 1483 591 1485 594
rect 1453 563 1455 573
rect 1483 563 1485 579
rect 1167 549 1169 558
rect 1085 528 1087 531
rect 1097 528 1099 531
rect 1128 528 1130 531
rect 1167 528 1169 545
rect 1175 542 1177 558
rect 1205 556 1207 559
rect 1324 546 1326 562
rect 1175 528 1177 538
rect 1205 528 1207 544
rect 1324 537 1326 540
rect 1358 535 1360 562
rect 1370 535 1372 562
rect 1401 529 1403 562
rect 1445 554 1447 557
rect 1453 554 1455 557
rect 1483 553 1485 557
rect 1167 519 1169 522
rect 1175 519 1177 522
rect 1205 518 1207 522
rect 1358 520 1360 523
rect 1370 520 1372 523
rect 1401 520 1403 523
rect 917 496 919 499
rect 929 496 931 499
rect 960 496 962 499
rect 1085 495 1087 498
rect 1097 495 1099 498
rect 1109 495 1111 498
rect 1139 495 1141 498
rect 805 487 807 490
rect 805 459 807 475
rect 839 466 841 493
rect 851 466 853 493
rect 882 460 884 493
rect 1358 488 1360 491
rect 1370 488 1372 491
rect 1401 488 1403 491
rect 923 470 925 473
rect 931 470 933 473
rect 805 450 807 453
rect 839 451 841 454
rect 851 451 853 454
rect 882 451 884 454
rect 1085 449 1087 483
rect 1097 449 1099 483
rect 1109 449 1111 483
rect 923 437 925 446
rect 805 427 807 430
rect 839 427 841 430
rect 851 427 853 430
rect 882 427 884 430
rect 923 416 925 433
rect 931 430 933 446
rect 961 444 963 447
rect 1139 446 1141 483
rect 1324 470 1326 473
rect 1184 464 1186 467
rect 1192 464 1194 467
rect 1200 464 1202 467
rect 1231 452 1233 455
rect 1324 442 1326 458
rect 1358 449 1360 476
rect 1370 449 1372 476
rect 1139 437 1141 440
rect 1085 434 1087 437
rect 1097 434 1099 437
rect 1109 434 1111 437
rect 931 416 933 426
rect 961 416 963 432
rect 1184 431 1186 440
rect 805 399 807 415
rect 805 390 807 393
rect 839 388 841 415
rect 851 388 853 415
rect 882 382 884 415
rect 923 407 925 410
rect 931 407 933 410
rect 961 406 963 410
rect 1184 403 1186 427
rect 1192 424 1194 440
rect 1192 403 1194 420
rect 1200 417 1202 440
rect 1231 424 1233 440
rect 1401 443 1403 476
rect 1445 453 1447 456
rect 1453 453 1455 456
rect 1324 433 1326 436
rect 1358 434 1360 437
rect 1370 434 1372 437
rect 1401 434 1403 437
rect 1445 420 1447 429
rect 1231 415 1233 418
rect 1200 403 1202 413
rect 1324 410 1326 413
rect 1358 410 1360 413
rect 1370 410 1372 413
rect 1401 410 1403 413
rect 1085 400 1087 403
rect 1097 400 1099 403
rect 1128 400 1130 403
rect 914 388 916 391
rect 926 388 928 391
rect 957 388 959 391
rect 1445 399 1447 416
rect 1453 413 1455 429
rect 1483 427 1485 430
rect 1453 399 1455 409
rect 1483 399 1485 415
rect 1184 394 1186 397
rect 1192 394 1194 397
rect 1200 394 1202 397
rect 839 373 841 376
rect 851 373 853 376
rect 882 373 884 376
rect 914 349 916 376
rect 926 349 928 376
rect 839 343 841 346
rect 851 343 853 346
rect 882 343 884 346
rect 957 343 959 376
rect 1085 361 1087 388
rect 1097 361 1099 388
rect 1128 355 1130 388
rect 1324 382 1326 398
rect 1324 373 1326 376
rect 1358 371 1360 398
rect 1370 371 1372 398
rect 1401 365 1403 398
rect 1445 390 1447 393
rect 1453 390 1455 393
rect 1483 389 1485 393
rect 1358 356 1360 359
rect 1370 356 1372 359
rect 1401 356 1403 359
rect 1085 346 1087 349
rect 1097 346 1099 349
rect 1128 346 1130 349
rect 914 334 916 337
rect 926 334 928 337
rect 957 334 959 337
rect 805 325 807 328
rect 805 297 807 313
rect 839 304 841 331
rect 851 304 853 331
rect 882 298 884 331
rect 1358 321 1360 324
rect 1370 321 1372 324
rect 1401 321 1403 324
rect 1085 311 1087 314
rect 1097 311 1099 314
rect 1109 311 1111 314
rect 1121 311 1123 314
rect 1146 311 1148 314
rect 926 308 928 311
rect 934 308 936 311
rect 805 288 807 291
rect 839 289 841 292
rect 851 289 853 292
rect 882 289 884 292
rect 1324 303 1326 306
rect 926 275 928 284
rect 805 265 807 268
rect 839 265 841 268
rect 851 265 853 268
rect 882 265 884 268
rect 926 254 928 271
rect 934 268 936 284
rect 964 282 966 285
rect 934 254 936 264
rect 964 254 966 270
rect 1085 258 1087 299
rect 1097 258 1099 299
rect 1109 258 1111 299
rect 1121 258 1123 299
rect 805 237 807 253
rect 805 228 807 231
rect 839 226 841 253
rect 851 226 853 253
rect 882 220 884 253
rect 926 245 928 248
rect 934 245 936 248
rect 964 244 966 248
rect 1146 255 1148 299
rect 1184 280 1186 283
rect 1192 280 1194 283
rect 1200 280 1202 283
rect 1208 280 1210 283
rect 1324 275 1326 291
rect 1358 282 1360 309
rect 1370 282 1372 309
rect 1401 276 1403 309
rect 1445 286 1447 289
rect 1453 286 1455 289
rect 1324 266 1326 269
rect 1358 267 1360 270
rect 1370 267 1372 270
rect 1401 267 1403 270
rect 1245 261 1247 264
rect 1146 246 1148 249
rect 1184 247 1186 256
rect 1085 243 1087 246
rect 1097 243 1099 246
rect 1109 243 1111 246
rect 1121 243 1123 246
rect 917 226 919 229
rect 929 226 931 229
rect 960 226 962 229
rect 839 211 841 214
rect 851 211 853 214
rect 882 211 884 214
rect 917 187 919 214
rect 929 187 931 214
rect 839 181 841 184
rect 851 181 853 184
rect 882 181 884 184
rect 960 181 962 214
rect 1085 213 1087 216
rect 1097 213 1099 216
rect 1109 213 1111 216
rect 1139 213 1141 216
rect 1184 211 1186 243
rect 1192 240 1194 256
rect 1192 211 1194 236
rect 1200 233 1202 256
rect 1200 211 1202 229
rect 1208 226 1210 256
rect 1445 253 1447 262
rect 1245 233 1247 249
rect 1324 243 1326 246
rect 1358 243 1360 246
rect 1370 243 1372 246
rect 1401 243 1403 246
rect 1445 232 1447 249
rect 1453 246 1455 262
rect 1483 260 1485 263
rect 1453 232 1455 242
rect 1483 232 1485 248
rect 1245 223 1247 227
rect 1208 211 1210 222
rect 1324 215 1326 231
rect 1324 206 1326 209
rect 1184 202 1186 205
rect 1192 202 1194 205
rect 1200 202 1202 205
rect 1208 202 1210 205
rect 1358 204 1360 231
rect 1370 204 1372 231
rect 917 172 919 175
rect 929 172 931 175
rect 960 172 962 175
rect 805 163 807 166
rect 805 135 807 151
rect 839 142 841 169
rect 851 142 853 169
rect 882 136 884 169
rect 1085 167 1087 201
rect 1097 167 1099 201
rect 1109 167 1111 201
rect 1139 164 1141 201
rect 1401 198 1403 231
rect 1445 223 1447 226
rect 1453 223 1455 226
rect 1483 222 1485 226
rect 1358 189 1360 192
rect 1370 189 1372 192
rect 1401 189 1403 192
rect 1139 155 1141 158
rect 1359 156 1361 159
rect 1371 156 1373 159
rect 1402 156 1404 159
rect 1085 152 1087 155
rect 1097 152 1099 155
rect 1109 152 1111 155
rect 923 146 925 149
rect 931 146 933 149
rect 805 126 807 129
rect 839 127 841 130
rect 851 127 853 130
rect 882 127 884 130
rect 1325 138 1327 141
rect 923 113 925 122
rect 805 103 807 106
rect 839 103 841 106
rect 851 103 853 106
rect 882 103 884 106
rect 923 92 925 109
rect 931 106 933 122
rect 961 120 963 123
rect 1085 120 1087 123
rect 1097 120 1099 123
rect 1128 120 1130 123
rect 1325 110 1327 126
rect 1359 117 1361 144
rect 1371 117 1373 144
rect 931 92 933 102
rect 961 92 963 108
rect 805 75 807 91
rect 805 66 807 69
rect 839 64 841 91
rect 851 64 853 91
rect 882 58 884 91
rect 923 83 925 86
rect 931 83 933 86
rect 961 82 963 86
rect 1085 81 1087 108
rect 1097 81 1099 108
rect 1128 75 1130 108
rect 1402 111 1404 144
rect 1446 121 1448 124
rect 1454 121 1456 124
rect 1325 101 1327 104
rect 1359 102 1361 105
rect 1371 102 1373 105
rect 1402 102 1404 105
rect 1446 88 1448 97
rect 1325 78 1327 81
rect 1359 78 1361 81
rect 1371 78 1373 81
rect 1402 78 1404 81
rect 914 64 916 67
rect 926 64 928 67
rect 957 64 959 67
rect 1085 66 1087 69
rect 1097 66 1099 69
rect 1128 66 1130 69
rect 1446 67 1448 84
rect 1454 81 1456 97
rect 1484 95 1486 98
rect 1454 67 1456 77
rect 1484 67 1486 83
rect 839 49 841 52
rect 851 49 853 52
rect 882 49 884 52
rect 914 25 916 52
rect 926 25 928 52
rect 957 19 959 52
rect 1325 50 1327 66
rect 1325 41 1327 44
rect 1359 39 1361 66
rect 1371 39 1373 66
rect 1402 33 1404 66
rect 1446 58 1448 61
rect 1454 58 1456 61
rect 1484 57 1486 61
rect 1359 24 1361 27
rect 1371 24 1373 27
rect 1402 24 1404 27
rect 914 10 916 13
rect 926 10 928 13
rect 957 10 959 13
<< polycontact >>
rect 835 640 839 644
rect 801 624 805 628
rect 847 637 851 641
rect 878 644 882 648
rect 1354 625 1358 629
rect 1320 609 1324 613
rect 924 595 928 599
rect 1366 622 1370 626
rect 1397 629 1401 633
rect 932 588 936 592
rect 960 581 964 585
rect 801 564 805 568
rect 835 560 839 564
rect 847 553 851 557
rect 878 564 882 568
rect 1081 553 1085 557
rect 1093 546 1097 550
rect 1124 557 1128 561
rect 913 521 917 525
rect 925 514 929 518
rect 956 525 960 529
rect 1443 580 1447 584
rect 1451 573 1455 577
rect 1479 566 1483 570
rect 1165 545 1169 549
rect 1320 549 1324 553
rect 1173 538 1177 542
rect 1201 531 1205 535
rect 1354 545 1358 549
rect 1366 538 1370 542
rect 1397 549 1401 553
rect 835 478 839 482
rect 801 462 805 466
rect 847 475 851 479
rect 878 482 882 486
rect 1081 466 1085 470
rect 1093 459 1097 463
rect 1105 452 1109 456
rect 1135 470 1139 474
rect 921 433 925 437
rect 1354 461 1358 465
rect 1320 445 1324 449
rect 1366 458 1370 462
rect 1397 465 1401 469
rect 929 426 933 430
rect 957 419 961 423
rect 1182 427 1186 431
rect 801 402 805 406
rect 835 398 839 402
rect 847 391 851 395
rect 878 402 882 406
rect 1190 420 1194 424
rect 1227 427 1231 431
rect 1198 413 1202 417
rect 1443 416 1447 420
rect 1451 409 1455 413
rect 1479 402 1483 406
rect 910 359 914 363
rect 922 352 926 356
rect 953 363 957 367
rect 1081 371 1085 375
rect 1093 364 1097 368
rect 1124 375 1128 379
rect 1320 385 1324 389
rect 1354 381 1358 385
rect 1366 374 1370 378
rect 1397 385 1401 389
rect 835 316 839 320
rect 801 300 805 304
rect 847 313 851 317
rect 878 320 882 324
rect 924 271 928 275
rect 1081 282 1085 286
rect 932 264 936 268
rect 960 257 964 261
rect 1093 275 1097 279
rect 1105 268 1109 272
rect 1117 261 1121 265
rect 1142 286 1146 290
rect 801 240 805 244
rect 835 236 839 240
rect 847 229 851 233
rect 878 240 882 244
rect 1354 294 1358 298
rect 1320 278 1324 282
rect 1366 291 1370 295
rect 1397 298 1401 302
rect 1182 243 1186 247
rect 913 197 917 201
rect 925 190 929 194
rect 956 201 960 205
rect 1190 236 1194 240
rect 1198 229 1202 233
rect 1443 249 1447 253
rect 1241 236 1245 240
rect 1451 242 1455 246
rect 1479 235 1483 239
rect 1206 222 1210 226
rect 1320 218 1324 222
rect 1354 214 1358 218
rect 1366 207 1370 211
rect 1397 218 1401 222
rect 1081 184 1085 188
rect 835 154 839 158
rect 801 138 805 142
rect 847 151 851 155
rect 878 158 882 162
rect 1093 177 1097 181
rect 1105 170 1109 174
rect 1135 188 1139 192
rect 1355 129 1359 133
rect 921 109 925 113
rect 1321 113 1325 117
rect 1367 126 1371 130
rect 1398 133 1402 137
rect 929 102 933 106
rect 957 95 961 99
rect 801 78 805 82
rect 835 74 839 78
rect 847 67 851 71
rect 878 78 882 82
rect 1081 91 1085 95
rect 1093 84 1097 88
rect 1124 95 1128 99
rect 1444 84 1448 88
rect 1452 77 1456 81
rect 1480 70 1484 74
rect 1321 53 1325 57
rect 910 35 914 39
rect 922 28 926 32
rect 953 39 957 43
rect 1355 49 1359 53
rect 1367 42 1371 46
rect 1398 53 1402 57
<< metal1 >>
rect 828 671 878 675
rect 834 667 838 671
rect 854 667 858 671
rect 794 653 818 657
rect 874 667 878 671
rect 1347 656 1397 660
rect 800 649 804 653
rect 844 648 848 655
rect 844 644 878 648
rect 888 646 892 655
rect 1353 652 1357 656
rect 1373 652 1377 656
rect 808 628 812 637
rect 822 640 835 644
rect 822 628 826 640
rect 843 635 847 641
rect 836 631 847 635
rect 856 628 860 644
rect 781 624 801 628
rect 808 624 826 628
rect 808 621 812 624
rect 888 642 910 646
rect 888 622 892 642
rect 800 611 804 615
rect 831 611 835 616
rect 874 611 878 616
rect 794 607 818 611
rect 828 607 878 611
rect 906 599 910 642
rect 913 636 952 640
rect 1313 638 1337 642
rect 1393 652 1397 656
rect 919 632 923 636
rect 948 614 952 636
rect 1319 634 1323 638
rect 1363 633 1367 640
rect 1363 629 1397 633
rect 1407 631 1411 640
rect 948 610 963 614
rect 1327 613 1331 622
rect 1341 625 1354 629
rect 1341 613 1345 625
rect 1362 620 1366 626
rect 1355 616 1366 620
rect 1375 613 1379 629
rect 794 593 818 597
rect 828 593 878 597
rect 906 595 924 599
rect 800 589 804 593
rect 834 589 838 593
rect 854 589 858 593
rect 874 589 878 593
rect 808 568 812 577
rect 844 568 848 577
rect 888 568 892 577
rect 906 588 932 592
rect 906 568 910 588
rect 939 585 943 608
rect 959 606 963 610
rect 1300 609 1320 613
rect 1327 609 1345 613
rect 1327 606 1331 609
rect 1407 627 1429 631
rect 1407 607 1411 627
rect 967 585 971 594
rect 1067 593 1286 597
rect 1319 596 1323 600
rect 1350 596 1354 601
rect 1393 596 1397 601
rect 1067 585 1071 593
rect 1074 586 1124 590
rect 1154 586 1193 590
rect 929 581 960 585
rect 967 581 1071 585
rect 1080 582 1084 586
rect 1100 582 1104 586
rect 929 578 933 581
rect 967 578 971 581
rect 919 568 923 572
rect 939 568 943 572
rect 959 568 963 572
rect 1120 582 1124 586
rect 1160 582 1164 586
rect 790 564 801 568
rect 808 564 830 568
rect 844 564 878 568
rect 888 564 910 568
rect 913 564 963 568
rect 808 561 812 564
rect 826 560 835 564
rect 800 551 804 555
rect 823 553 847 557
rect 794 547 818 551
rect 785 527 789 546
rect 823 536 827 553
rect 856 550 860 564
rect 888 544 892 564
rect 1090 561 1094 570
rect 1134 561 1138 570
rect 906 554 956 558
rect 1090 557 1124 561
rect 1134 557 1151 561
rect 1189 564 1193 586
rect 1189 560 1204 564
rect 912 550 916 554
rect 932 550 936 554
rect 952 550 956 554
rect 1026 553 1081 557
rect 831 533 835 538
rect 874 533 878 538
rect 828 530 878 533
rect 922 529 926 538
rect 966 529 970 538
rect 1026 529 1030 553
rect 785 525 893 527
rect 922 525 956 529
rect 966 525 1030 529
rect 785 523 913 525
rect 889 521 913 523
rect 781 518 886 520
rect 781 516 925 518
rect 882 514 925 516
rect 828 509 878 513
rect 934 511 938 525
rect 834 505 838 509
rect 854 505 858 509
rect 794 491 818 495
rect 874 505 878 509
rect 966 505 970 525
rect 909 494 913 499
rect 952 494 956 499
rect 800 487 804 491
rect 844 486 848 493
rect 844 482 878 486
rect 888 484 892 493
rect 906 490 956 494
rect 808 466 812 475
rect 822 478 835 482
rect 822 466 826 478
rect 843 473 847 479
rect 836 469 847 473
rect 856 466 860 482
rect 781 462 801 466
rect 808 462 826 466
rect 808 459 812 462
rect 888 480 907 484
rect 888 460 892 480
rect 800 449 804 453
rect 831 449 835 454
rect 874 449 878 454
rect 794 445 818 449
rect 828 445 878 449
rect 903 437 907 480
rect 910 474 949 478
rect 916 470 920 474
rect 945 452 949 474
rect 1026 456 1030 525
rect 1043 546 1093 550
rect 1043 466 1047 546
rect 1102 543 1106 557
rect 1134 537 1138 557
rect 1147 549 1151 557
rect 1147 545 1165 549
rect 1147 538 1173 542
rect 1077 526 1081 531
rect 1120 526 1124 531
rect 1074 522 1124 526
rect 1147 519 1151 538
rect 1180 535 1184 558
rect 1200 556 1204 560
rect 1208 535 1212 544
rect 1282 544 1286 593
rect 1313 592 1337 596
rect 1347 592 1397 596
rect 1425 584 1429 627
rect 1432 621 1471 625
rect 1438 617 1442 621
rect 1467 599 1471 621
rect 1467 595 1482 599
rect 1313 578 1337 582
rect 1347 578 1397 582
rect 1425 580 1443 584
rect 1319 574 1323 578
rect 1353 574 1357 578
rect 1373 574 1377 578
rect 1393 574 1397 578
rect 1327 553 1331 562
rect 1363 553 1367 562
rect 1407 553 1411 562
rect 1425 573 1451 577
rect 1425 553 1429 573
rect 1458 570 1462 593
rect 1478 591 1482 595
rect 1486 570 1490 579
rect 1448 566 1479 570
rect 1486 566 1494 570
rect 1448 563 1452 566
rect 1486 563 1490 566
rect 1438 553 1442 557
rect 1458 553 1462 557
rect 1478 553 1482 557
rect 1309 549 1320 553
rect 1327 549 1349 553
rect 1363 549 1397 553
rect 1407 549 1429 553
rect 1432 549 1482 553
rect 1313 544 1316 549
rect 1327 546 1331 549
rect 1282 540 1316 544
rect 1345 545 1354 549
rect 1319 536 1323 540
rect 1342 538 1366 542
rect 1170 531 1201 535
rect 1208 531 1284 535
rect 1313 532 1337 536
rect 1170 528 1174 531
rect 1208 528 1212 531
rect 1051 515 1151 519
rect 1160 518 1164 522
rect 1180 518 1184 522
rect 1200 518 1204 522
rect 1051 475 1055 515
rect 1154 514 1204 518
rect 1074 499 1135 503
rect 1080 495 1084 499
rect 1102 495 1106 499
rect 1131 495 1135 499
rect 1090 474 1094 483
rect 1112 474 1116 483
rect 1145 474 1149 483
rect 1090 470 1135 474
rect 1145 470 1168 474
rect 1048 463 1061 466
rect 1048 462 1093 463
rect 1057 459 1093 462
rect 1026 452 1105 456
rect 945 448 960 452
rect 794 431 818 435
rect 828 431 878 435
rect 903 433 921 437
rect 800 427 804 431
rect 834 427 838 431
rect 854 427 858 431
rect 874 427 878 431
rect 808 406 812 415
rect 844 406 848 415
rect 888 406 892 415
rect 903 426 929 430
rect 903 406 907 426
rect 936 423 940 446
rect 956 444 960 448
rect 964 423 968 432
rect 926 419 957 423
rect 964 419 1017 423
rect 926 416 930 419
rect 964 416 968 419
rect 916 406 920 410
rect 936 406 940 410
rect 956 406 960 410
rect 790 402 801 406
rect 808 402 830 406
rect 844 402 878 406
rect 888 402 907 406
rect 910 402 960 406
rect 808 399 812 402
rect 826 398 835 402
rect 800 389 804 393
rect 823 391 847 395
rect 794 385 818 389
rect 785 365 789 384
rect 823 374 827 391
rect 856 388 860 402
rect 888 382 892 402
rect 903 392 953 396
rect 909 388 913 392
rect 929 388 933 392
rect 949 388 953 392
rect 831 371 835 376
rect 874 371 878 376
rect 828 368 878 371
rect 919 367 923 376
rect 963 367 967 376
rect 785 363 893 365
rect 919 363 953 367
rect 963 363 1016 367
rect 785 361 910 363
rect 889 359 910 361
rect 781 356 886 358
rect 781 354 922 356
rect 882 352 922 354
rect 828 347 878 351
rect 931 349 935 363
rect 834 343 838 347
rect 854 343 858 347
rect 794 329 818 333
rect 874 343 878 347
rect 963 343 967 363
rect 906 332 910 337
rect 949 332 953 337
rect 800 325 804 329
rect 844 324 848 331
rect 844 320 878 324
rect 888 322 892 331
rect 903 328 953 332
rect 808 304 812 313
rect 822 316 835 320
rect 822 304 826 316
rect 843 311 847 317
rect 836 307 847 311
rect 856 304 860 320
rect 781 300 801 304
rect 808 300 826 304
rect 808 297 812 300
rect 888 318 910 322
rect 888 298 892 318
rect 800 287 804 291
rect 831 287 835 292
rect 874 287 878 292
rect 794 283 818 287
rect 828 283 878 287
rect 906 275 910 318
rect 913 312 952 316
rect 919 308 923 312
rect 948 290 952 312
rect 948 286 963 290
rect 794 269 818 273
rect 828 269 878 273
rect 906 271 924 275
rect 800 265 804 269
rect 834 265 838 269
rect 854 265 858 269
rect 874 265 878 269
rect 808 244 812 253
rect 844 244 848 253
rect 888 244 892 253
rect 906 264 932 268
rect 906 244 910 264
rect 939 261 943 284
rect 959 282 963 286
rect 1026 265 1030 452
rect 1112 449 1116 470
rect 1043 423 1047 442
rect 1039 419 1047 423
rect 1043 272 1047 419
rect 1052 368 1056 443
rect 1145 446 1149 470
rect 1077 432 1081 437
rect 1131 432 1135 440
rect 1074 428 1135 432
rect 1164 431 1168 470
rect 1171 468 1216 472
rect 1177 464 1181 468
rect 1212 460 1216 468
rect 1212 456 1230 460
rect 1226 452 1230 456
rect 1205 431 1209 440
rect 1234 431 1238 440
rect 1164 427 1182 431
rect 1205 427 1227 431
rect 1234 427 1277 431
rect 1147 420 1190 424
rect 1074 404 1124 408
rect 1080 400 1084 404
rect 1100 400 1104 404
rect 1120 400 1124 404
rect 1090 379 1094 388
rect 1134 379 1138 388
rect 1147 379 1151 420
rect 1060 368 1064 376
rect 1090 375 1124 379
rect 1134 375 1151 379
rect 1163 413 1198 417
rect 1052 364 1093 368
rect 1052 285 1056 364
rect 1102 361 1106 375
rect 1134 355 1138 375
rect 1077 344 1081 349
rect 1120 344 1124 349
rect 1074 340 1124 344
rect 1163 337 1167 413
rect 1205 410 1209 427
rect 1234 424 1238 427
rect 1226 414 1230 418
rect 1187 406 1209 410
rect 1187 403 1191 406
rect 1205 403 1209 406
rect 1212 410 1230 414
rect 1177 393 1181 397
rect 1195 393 1199 397
rect 1212 393 1216 410
rect 1171 389 1216 393
rect 1060 333 1167 337
rect 1060 302 1064 333
rect 1074 315 1142 319
rect 1080 311 1084 315
rect 1102 311 1106 315
rect 1124 311 1128 315
rect 1138 311 1142 315
rect 1090 290 1094 299
rect 1114 290 1118 299
rect 1152 290 1156 299
rect 1090 286 1142 290
rect 1152 286 1168 290
rect 1061 282 1081 286
rect 1043 268 1105 272
rect 1026 261 1117 265
rect 929 257 960 261
rect 1124 258 1128 286
rect 929 254 933 257
rect 919 244 923 248
rect 939 244 943 248
rect 959 244 963 248
rect 790 240 801 244
rect 808 240 830 244
rect 844 240 878 244
rect 888 240 910 244
rect 913 240 963 244
rect 808 237 812 240
rect 826 236 835 240
rect 800 227 804 231
rect 823 229 847 233
rect 794 223 818 227
rect 785 203 789 222
rect 823 212 827 229
rect 856 226 860 240
rect 888 220 892 240
rect 906 230 956 234
rect 912 226 916 230
rect 932 226 936 230
rect 952 226 956 230
rect 831 209 835 214
rect 874 209 878 214
rect 828 206 878 209
rect 922 205 926 214
rect 966 205 970 214
rect 1039 205 1043 252
rect 785 201 893 203
rect 922 201 956 205
rect 966 201 1043 205
rect 785 199 913 201
rect 889 197 913 199
rect 781 194 886 196
rect 781 192 925 194
rect 882 190 925 192
rect 828 185 878 189
rect 934 187 938 201
rect 834 181 838 185
rect 854 181 858 185
rect 794 167 818 171
rect 874 181 878 185
rect 966 181 970 201
rect 909 170 913 175
rect 952 170 956 175
rect 800 163 804 167
rect 844 162 848 169
rect 844 158 878 162
rect 888 160 892 169
rect 906 166 956 170
rect 808 142 812 151
rect 822 154 835 158
rect 822 142 826 154
rect 843 149 847 155
rect 836 145 847 149
rect 856 142 860 158
rect 781 138 801 142
rect 808 138 826 142
rect 808 135 812 138
rect 888 156 907 160
rect 888 136 892 156
rect 800 125 804 129
rect 831 125 835 130
rect 874 125 878 130
rect 794 121 818 125
rect 828 121 878 125
rect 903 113 907 156
rect 910 150 949 154
rect 916 146 920 150
rect 945 128 949 150
rect 945 124 960 128
rect 794 107 818 111
rect 828 107 878 111
rect 903 109 921 113
rect 800 103 804 107
rect 834 103 838 107
rect 854 103 858 107
rect 874 103 878 107
rect 808 82 812 91
rect 844 82 848 91
rect 888 82 892 91
rect 903 102 929 106
rect 903 82 907 102
rect 936 99 940 122
rect 956 120 960 124
rect 964 99 968 108
rect 926 95 957 99
rect 964 95 1030 99
rect 926 92 930 95
rect 964 92 968 95
rect 916 82 920 86
rect 936 82 940 86
rect 1039 88 1043 201
rect 1051 174 1055 252
rect 1060 188 1064 252
rect 1152 255 1156 286
rect 1077 241 1081 246
rect 1138 241 1142 249
rect 1164 247 1168 286
rect 1171 284 1225 288
rect 1177 280 1181 284
rect 1221 269 1225 284
rect 1221 265 1244 269
rect 1164 243 1182 247
rect 1074 237 1142 241
rect 1213 240 1217 256
rect 1240 261 1244 265
rect 1248 240 1252 249
rect 1157 236 1190 240
rect 1213 236 1241 240
rect 1248 236 1256 240
rect 1074 217 1135 221
rect 1080 213 1084 217
rect 1102 213 1106 217
rect 1131 213 1135 217
rect 1090 192 1094 201
rect 1112 192 1116 201
rect 1145 192 1149 201
rect 1157 192 1161 236
rect 1090 188 1135 192
rect 1145 188 1161 192
rect 1164 222 1206 226
rect 1060 184 1081 188
rect 1060 183 1064 184
rect 1051 170 1105 174
rect 1112 167 1116 188
rect 1059 99 1063 161
rect 1145 164 1149 188
rect 1077 150 1081 155
rect 1131 150 1135 158
rect 1074 146 1135 150
rect 1074 124 1124 128
rect 1080 120 1084 124
rect 1100 120 1104 124
rect 1120 120 1124 124
rect 1052 95 1063 99
rect 1090 99 1094 108
rect 1134 99 1138 108
rect 1164 99 1168 222
rect 1213 218 1217 236
rect 1248 233 1252 236
rect 1240 223 1244 227
rect 1187 214 1217 218
rect 1226 219 1244 223
rect 1187 211 1191 214
rect 1203 211 1207 214
rect 1177 201 1181 205
rect 1195 201 1199 205
rect 1213 201 1217 205
rect 1226 201 1230 219
rect 1171 197 1230 201
rect 1273 125 1277 427
rect 1280 290 1284 531
rect 1342 521 1346 538
rect 1375 535 1379 549
rect 1407 529 1411 549
rect 1350 518 1354 523
rect 1393 518 1397 523
rect 1347 514 1397 518
rect 1347 492 1397 496
rect 1353 488 1357 492
rect 1373 488 1377 492
rect 1313 474 1337 478
rect 1393 488 1397 492
rect 1319 470 1323 474
rect 1363 469 1367 476
rect 1363 465 1397 469
rect 1407 467 1411 476
rect 1327 449 1331 458
rect 1341 461 1354 465
rect 1341 449 1345 461
rect 1362 456 1366 462
rect 1355 452 1366 456
rect 1375 449 1379 465
rect 1300 445 1320 449
rect 1327 445 1345 449
rect 1327 442 1331 445
rect 1407 463 1429 467
rect 1407 443 1411 463
rect 1319 432 1323 436
rect 1350 432 1354 437
rect 1393 432 1397 437
rect 1313 428 1337 432
rect 1347 428 1397 432
rect 1425 420 1429 463
rect 1432 457 1471 461
rect 1438 453 1442 457
rect 1467 435 1471 457
rect 1467 431 1482 435
rect 1313 414 1337 418
rect 1347 414 1397 418
rect 1425 416 1443 420
rect 1319 410 1323 414
rect 1353 410 1357 414
rect 1373 410 1377 414
rect 1393 410 1397 414
rect 1327 389 1331 398
rect 1363 389 1367 398
rect 1407 389 1411 398
rect 1425 409 1451 413
rect 1425 389 1429 409
rect 1458 406 1462 429
rect 1478 427 1482 431
rect 1486 406 1490 415
rect 1448 402 1479 406
rect 1486 402 1494 406
rect 1448 399 1452 402
rect 1486 399 1490 402
rect 1438 389 1442 393
rect 1458 389 1462 393
rect 1478 389 1482 393
rect 1309 385 1320 389
rect 1327 385 1349 389
rect 1363 385 1397 389
rect 1407 385 1429 389
rect 1432 385 1482 389
rect 1327 382 1331 385
rect 1345 381 1354 385
rect 1319 372 1323 376
rect 1342 374 1366 378
rect 1313 368 1337 372
rect 1342 357 1346 374
rect 1375 371 1379 385
rect 1407 365 1411 385
rect 1350 354 1354 359
rect 1393 354 1397 359
rect 1347 351 1397 354
rect 1347 325 1397 329
rect 1353 321 1357 325
rect 1373 321 1377 325
rect 1313 307 1337 311
rect 1393 321 1397 325
rect 1319 303 1323 307
rect 1363 302 1367 309
rect 1363 298 1397 302
rect 1407 300 1411 309
rect 1280 286 1313 290
rect 1309 282 1313 286
rect 1327 282 1331 291
rect 1341 294 1354 298
rect 1341 282 1345 294
rect 1362 289 1366 295
rect 1355 285 1366 289
rect 1375 282 1379 298
rect 1300 278 1320 282
rect 1327 278 1345 282
rect 1327 275 1331 278
rect 1407 296 1429 300
rect 1407 276 1411 296
rect 1319 265 1323 269
rect 1350 265 1354 270
rect 1393 265 1397 270
rect 1313 261 1337 265
rect 1347 261 1397 265
rect 1425 253 1429 296
rect 1432 290 1471 294
rect 1438 286 1442 290
rect 1467 268 1471 290
rect 1467 264 1482 268
rect 1313 247 1337 251
rect 1347 247 1397 251
rect 1425 249 1443 253
rect 1319 243 1323 247
rect 1353 243 1357 247
rect 1373 243 1377 247
rect 1393 243 1397 247
rect 1327 222 1331 231
rect 1363 222 1367 231
rect 1407 222 1411 231
rect 1425 242 1451 246
rect 1425 222 1429 242
rect 1458 239 1462 262
rect 1478 260 1482 264
rect 1486 239 1490 248
rect 1448 235 1479 239
rect 1486 235 1494 239
rect 1448 232 1452 235
rect 1486 232 1490 235
rect 1438 222 1442 226
rect 1458 222 1462 226
rect 1478 222 1482 226
rect 1309 218 1320 222
rect 1327 218 1349 222
rect 1363 218 1397 222
rect 1407 218 1429 222
rect 1432 218 1482 222
rect 1327 215 1331 218
rect 1345 214 1354 218
rect 1319 205 1323 209
rect 1342 207 1366 211
rect 1313 201 1337 205
rect 1342 190 1346 207
rect 1375 204 1379 218
rect 1407 198 1411 218
rect 1350 187 1354 192
rect 1393 187 1397 192
rect 1347 184 1397 187
rect 1348 160 1398 164
rect 1354 156 1358 160
rect 1374 156 1378 160
rect 1314 142 1338 146
rect 1394 156 1398 160
rect 1320 138 1324 142
rect 1364 137 1368 144
rect 1364 133 1398 137
rect 1408 135 1412 144
rect 1273 121 1314 125
rect 1310 117 1314 121
rect 1328 117 1332 126
rect 1342 129 1355 133
rect 1342 117 1346 129
rect 1363 124 1367 130
rect 1356 120 1367 124
rect 1376 117 1380 133
rect 1301 113 1321 117
rect 1328 113 1346 117
rect 1328 110 1332 113
rect 1408 131 1430 135
rect 1408 111 1412 131
rect 1320 100 1324 104
rect 1351 100 1355 105
rect 1394 100 1398 105
rect 1090 95 1124 99
rect 1134 95 1168 99
rect 1314 96 1338 100
rect 1348 96 1398 100
rect 1059 91 1081 95
rect 956 82 960 86
rect 1039 84 1093 88
rect 790 78 801 82
rect 808 78 830 82
rect 844 78 878 82
rect 888 78 907 82
rect 910 78 960 82
rect 1102 81 1106 95
rect 808 75 812 78
rect 826 74 835 78
rect 800 65 804 69
rect 823 67 847 71
rect 794 61 818 65
rect 785 41 789 60
rect 823 50 827 67
rect 856 64 860 78
rect 888 58 892 78
rect 903 68 953 72
rect 909 64 913 68
rect 929 64 933 68
rect 949 64 953 68
rect 1134 75 1138 95
rect 1426 88 1430 131
rect 1433 125 1472 129
rect 1439 121 1443 125
rect 1468 103 1472 125
rect 1468 99 1483 103
rect 1314 82 1338 86
rect 1348 82 1398 86
rect 1426 84 1444 88
rect 1320 78 1324 82
rect 1354 78 1358 82
rect 1374 78 1378 82
rect 1077 64 1081 69
rect 1120 64 1124 69
rect 1394 78 1398 82
rect 1074 60 1124 64
rect 1328 57 1332 66
rect 1364 57 1368 66
rect 1408 57 1412 66
rect 1426 77 1452 81
rect 1426 57 1430 77
rect 1459 74 1463 97
rect 1479 95 1483 99
rect 1487 74 1491 83
rect 1449 70 1480 74
rect 1487 70 1495 74
rect 1449 67 1453 70
rect 1487 67 1491 70
rect 1439 57 1443 61
rect 1459 57 1463 61
rect 1479 57 1483 61
rect 1310 53 1321 57
rect 1328 53 1350 57
rect 1364 53 1398 57
rect 1408 53 1430 57
rect 1433 53 1483 57
rect 831 47 835 52
rect 874 47 878 52
rect 828 44 878 47
rect 919 43 923 52
rect 1328 50 1332 53
rect 1346 49 1355 53
rect 785 39 893 41
rect 919 39 953 43
rect 1320 40 1324 44
rect 1343 42 1367 46
rect 785 37 910 39
rect 889 35 910 37
rect 781 32 886 34
rect 781 30 922 32
rect 882 28 922 30
rect 931 25 935 39
rect 1314 36 1338 40
rect 1343 25 1347 42
rect 1376 39 1380 53
rect 1408 33 1412 53
rect 1351 22 1355 27
rect 1394 22 1398 27
rect 1348 18 1398 22
rect 906 8 910 13
rect 949 8 953 13
rect 903 4 953 8
<< m2contact >>
rect 831 631 836 636
rect 776 623 781 628
rect 1350 616 1355 621
rect 1295 608 1300 613
rect 785 563 790 568
rect 785 546 790 551
rect 818 536 823 541
rect 776 516 781 521
rect 831 469 836 474
rect 776 461 781 466
rect 1038 518 1043 523
rect 1030 501 1035 506
rect 1304 548 1309 553
rect 1051 470 1056 475
rect 1043 461 1048 466
rect 1017 419 1022 424
rect 785 401 790 406
rect 785 384 790 389
rect 818 374 823 379
rect 1016 363 1021 368
rect 776 354 781 359
rect 831 307 836 312
rect 776 299 781 304
rect 1043 442 1048 447
rect 1052 443 1057 448
rect 1034 419 1039 424
rect 1060 376 1065 381
rect 1060 297 1065 302
rect 1051 280 1056 285
rect 1060 277 1065 282
rect 1039 252 1044 257
rect 1050 252 1055 257
rect 785 239 790 244
rect 785 222 790 227
rect 818 212 823 217
rect 776 192 781 197
rect 831 145 836 150
rect 776 137 781 142
rect 1030 95 1035 100
rect 1060 252 1065 257
rect 1059 178 1064 183
rect 1059 161 1064 166
rect 1047 95 1052 100
rect 1063 136 1068 141
rect 1337 521 1342 526
rect 1350 452 1355 457
rect 1295 444 1300 449
rect 1304 384 1309 389
rect 1337 357 1342 362
rect 1350 285 1355 290
rect 1295 277 1300 282
rect 1304 217 1309 222
rect 1337 190 1342 195
rect 1351 120 1356 125
rect 1296 112 1301 117
rect 785 77 790 82
rect 785 60 790 65
rect 818 50 823 55
rect 1305 52 1310 57
rect 776 30 781 35
rect 1338 25 1343 30
<< metal2 >>
rect 785 660 825 664
rect 776 540 780 623
rect 785 568 789 660
rect 821 648 825 660
rect 821 645 831 648
rect 827 631 831 645
rect 1304 645 1344 649
rect 785 551 789 563
rect 776 536 818 540
rect 776 521 780 536
rect 1295 525 1299 608
rect 1304 553 1308 645
rect 1340 633 1344 645
rect 1340 630 1350 633
rect 1346 616 1350 630
rect 1295 521 1337 525
rect 1038 514 1041 518
rect 1038 510 1327 514
rect 785 498 825 502
rect 1035 502 1291 506
rect 776 378 780 461
rect 785 406 789 498
rect 821 486 825 498
rect 821 483 831 486
rect 827 469 831 483
rect 1043 447 1047 461
rect 1052 448 1056 470
rect 1072 466 1081 470
rect 1022 419 1034 423
rect 785 389 789 401
rect 776 374 818 378
rect 1039 376 1060 380
rect 776 359 780 374
rect 1039 367 1043 376
rect 1021 363 1043 367
rect 1072 375 1076 466
rect 1287 440 1291 502
rect 1323 485 1327 510
rect 1304 481 1344 485
rect 1295 440 1299 444
rect 1287 436 1299 440
rect 1072 371 1081 375
rect 785 336 825 340
rect 776 216 780 299
rect 785 244 789 336
rect 821 324 825 336
rect 1072 324 1076 371
rect 1295 361 1299 436
rect 1304 389 1308 481
rect 1340 469 1344 481
rect 1340 466 1350 469
rect 1346 452 1350 466
rect 1295 357 1337 361
rect 821 321 831 324
rect 827 307 831 321
rect 1072 320 1308 324
rect 1060 293 1064 297
rect 1039 289 1064 293
rect 967 261 971 270
rect 967 257 1035 261
rect 967 254 971 257
rect 1031 248 1035 257
rect 1039 257 1043 289
rect 1051 257 1055 280
rect 1061 257 1065 277
rect 1072 279 1076 320
rect 1304 318 1308 320
rect 1304 314 1344 318
rect 1072 275 1093 279
rect 1072 248 1076 275
rect 1031 244 1076 248
rect 785 227 789 239
rect 974 229 1030 233
rect 776 212 818 216
rect 776 197 780 212
rect 785 174 825 178
rect 776 54 780 137
rect 785 82 789 174
rect 821 162 825 174
rect 821 159 831 162
rect 827 145 831 159
rect 785 65 789 77
rect 776 50 818 54
rect 776 35 780 50
rect 963 43 967 52
rect 974 43 978 229
rect 1072 181 1076 244
rect 1089 229 1198 233
rect 1295 194 1299 277
rect 1304 222 1308 314
rect 1340 302 1344 314
rect 1340 299 1350 302
rect 1346 285 1350 299
rect 1295 190 1337 194
rect 1059 166 1063 178
rect 1072 177 1093 181
rect 1305 149 1345 153
rect 1305 141 1309 149
rect 1068 137 1309 141
rect 1035 95 1047 99
rect 963 39 978 43
rect 963 19 967 39
rect 1296 29 1300 112
rect 1305 57 1309 137
rect 1341 137 1345 149
rect 1341 134 1351 137
rect 1347 120 1351 134
rect 1296 25 1338 29
<< m3contact >>
rect 1030 228 1035 233
rect 1084 228 1089 233
<< metal3 >>
rect 1035 229 1084 233
<< labels >>
rlabel metal1 1321 639 1321 639 5 VDD
rlabel metal1 1324 594 1324 594 1 GND
rlabel metal1 1321 579 1321 579 5 VDD
rlabel metal1 1324 534 1324 534 1 GND
rlabel metal1 1365 580 1365 580 5 VDD
rlabel metal1 1379 516 1379 516 1 GND
rlabel metal1 1365 658 1365 658 5 VDD
rlabel metal1 1379 594 1379 594 1 GND
rlabel metal1 1449 623 1449 623 5 VDD
rlabel metal1 1450 551 1450 551 1 GND
rlabel ndcontact 1321 603 1321 603 1 GND
rlabel pdcontact 1321 628 1321 628 1 VDD
rlabel ndcontact 1352 607 1352 607 1 GND
rlabel pdcontact 1355 646 1355 646 1 VDD
rlabel pdcontact 1375 646 1375 646 1 VDD
rlabel pdcontact 1395 646 1395 646 1 VDD
rlabel ndcontact 1395 604 1395 604 1 GND
rlabel ndcontact 1440 560 1440 560 1 GND
rlabel ndcontact 1460 560 1460 560 1 GND
rlabel ndcontact 1480 560 1480 560 1 GND
rlabel pdcontact 1480 585 1480 585 1 VDD
rlabel pdcontact 1480 254 1480 254 1 VDD
rlabel ndcontact 1480 229 1480 229 1 GND
rlabel ndcontact 1460 229 1460 229 1 GND
rlabel ndcontact 1440 229 1440 229 1 GND
rlabel ndcontact 1395 195 1395 195 1 GND
rlabel pdcontact 1395 237 1395 237 1 VDD
rlabel ndcontact 1395 273 1395 273 1 GND
rlabel pdcontact 1395 315 1395 315 1 VDD
rlabel pdcontact 1375 315 1375 315 1 VDD
rlabel pdcontact 1355 315 1355 315 1 VDD
rlabel ndcontact 1352 276 1352 276 1 GND
rlabel pdcontact 1375 237 1375 237 1 VDD
rlabel pdcontact 1355 237 1355 237 1 VDD
rlabel ndcontact 1352 198 1352 198 1 GND
rlabel pdcontact 1321 297 1321 297 1 VDD
rlabel ndcontact 1321 272 1321 272 1 GND
rlabel pdcontact 1321 237 1321 237 1 VDD
rlabel ndcontact 1321 212 1321 212 1 GND
rlabel metal1 1450 220 1450 220 1 GND
rlabel metal1 1449 292 1449 292 5 VDD
rlabel metal1 1379 263 1379 263 1 GND
rlabel metal1 1365 327 1365 327 5 VDD
rlabel metal1 1379 185 1379 185 1 GND
rlabel metal1 1365 249 1365 249 5 VDD
rlabel metal1 1324 203 1324 203 1 GND
rlabel metal1 1321 248 1321 248 5 VDD
rlabel metal1 1324 263 1324 263 1 GND
rlabel metal1 1321 308 1321 308 5 VDD
rlabel metal1 1321 475 1321 475 5 VDD
rlabel metal1 1324 430 1324 430 1 GND
rlabel metal1 1321 415 1321 415 5 VDD
rlabel metal1 1324 370 1324 370 1 GND
rlabel metal1 1365 416 1365 416 5 VDD
rlabel metal1 1379 352 1379 352 1 GND
rlabel metal1 1365 494 1365 494 5 VDD
rlabel metal1 1379 430 1379 430 1 GND
rlabel metal1 1449 459 1449 459 5 VDD
rlabel metal1 1450 387 1450 387 1 GND
rlabel ndcontact 1321 379 1321 379 1 GND
rlabel pdcontact 1321 404 1321 404 1 VDD
rlabel ndcontact 1321 439 1321 439 1 GND
rlabel pdcontact 1321 464 1321 464 1 VDD
rlabel ndcontact 1352 365 1352 365 1 GND
rlabel pdcontact 1355 404 1355 404 1 VDD
rlabel pdcontact 1375 404 1375 404 1 VDD
rlabel ndcontact 1352 443 1352 443 1 GND
rlabel pdcontact 1355 482 1355 482 1 VDD
rlabel pdcontact 1375 482 1375 482 1 VDD
rlabel pdcontact 1395 482 1395 482 1 VDD
rlabel ndcontact 1395 440 1395 440 1 GND
rlabel pdcontact 1395 404 1395 404 1 VDD
rlabel ndcontact 1395 362 1395 362 1 GND
rlabel ndcontact 1440 396 1440 396 1 GND
rlabel ndcontact 1460 396 1460 396 1 GND
rlabel ndcontact 1480 396 1480 396 1 GND
rlabel pdcontact 1480 421 1480 421 1 VDD
rlabel metal1 1322 143 1322 143 5 VDD
rlabel metal1 1325 98 1325 98 1 GND
rlabel metal1 1322 83 1322 83 5 VDD
rlabel metal1 1325 38 1325 38 1 GND
rlabel metal1 1366 84 1366 84 5 VDD
rlabel metal1 1380 20 1380 20 1 GND
rlabel metal1 1366 162 1366 162 5 VDD
rlabel metal1 1380 98 1380 98 1 GND
rlabel metal1 1450 127 1450 127 5 VDD
rlabel metal1 1451 55 1451 55 1 GND
rlabel ndcontact 1322 47 1322 47 1 GND
rlabel pdcontact 1322 72 1322 72 1 VDD
rlabel ndcontact 1322 107 1322 107 1 GND
rlabel pdcontact 1322 132 1322 132 1 VDD
rlabel ndcontact 1353 33 1353 33 1 GND
rlabel pdcontact 1356 72 1356 72 1 VDD
rlabel pdcontact 1376 72 1376 72 1 VDD
rlabel ndcontact 1353 111 1353 111 1 GND
rlabel pdcontact 1356 150 1356 150 1 VDD
rlabel pdcontact 1376 150 1376 150 1 VDD
rlabel pdcontact 1396 150 1396 150 1 VDD
rlabel ndcontact 1396 108 1396 108 1 GND
rlabel pdcontact 1396 72 1396 72 1 VDD
rlabel ndcontact 1396 30 1396 30 1 GND
rlabel ndcontact 1441 64 1441 64 1 GND
rlabel ndcontact 1461 64 1461 64 1 GND
rlabel ndcontact 1481 64 1481 64 1 GND
rlabel pdcontact 1481 89 1481 89 1 VDD
rlabel polycontact 1322 551 1322 551 1 p0
rlabel pdcontact 1329 568 1329 568 1 p0_bar
rlabel polycontact 1356 547 1356 547 1 p0_bar
rlabel polycontact 1368 540 1368 540 1 c0
rlabel polycontact 1322 611 1322 611 1 c0
rlabel pdcontact 1329 628 1329 628 1 c0_bar
rlabel polycontact 1356 627 1356 627 1 c0_bar
rlabel polycontact 1368 624 1368 624 1 p0
rlabel metal1 1492 568 1492 568 7 s0
rlabel ndcontact 1488 560 1488 560 1 s0
rlabel pdcontact 1488 585 1488 585 1 s0
rlabel pdcontact 1440 605 1440 605 1 vdd
rlabel pdcontact 1365 646 1365 646 1 a1n
rlabel ndiffusion 1365 607 1365 607 1 a1m
rlabel ndcontact 1377 607 1377 607 1 a1n
rlabel polycontact 1399 631 1399 631 1 a1n
rlabel ndcontact 1409 604 1409 604 1 outa1
rlabel pdcontact 1409 646 1409 646 1 outa1
rlabel polycontact 1445 582 1445 582 1 outa1
rlabel polycontact 1453 575 1453 575 1 outa2
rlabel polycontact 1481 568 1481 568 1 s0_bar
rlabel ndcontact 1450 560 1450 560 1 s0_bar
rlabel pdcontact 1460 605 1460 605 1 s0_bar
rlabel pdcontact 1409 568 1409 568 1 outa2
rlabel ndcontact 1409 526 1409 526 1 outa2
rlabel polycontact 1399 551 1399 551 1 a2n
rlabel pdcontact 1365 568 1365 568 1 a2n
rlabel ndcontact 1377 529 1377 529 1 a2n
rlabel ndiffusion 1365 529 1365 529 1 a2m
rlabel polycontact 1322 387 1322 387 1 p1
rlabel ndcontact 1329 379 1329 379 1 p1_bar
rlabel pdcontact 1329 404 1329 404 1 p1_bar
rlabel polycontact 1356 383 1356 383 1 p1_bar
rlabel pdcontact 1365 404 1365 404 1 b2n
rlabel ndcontact 1377 365 1377 365 1 b2n
rlabel ndiffusion 1365 365 1365 365 1 b2m
rlabel polycontact 1399 387 1399 387 1 b2n
rlabel pdcontact 1409 404 1409 404 1 outb2
rlabel ndcontact 1409 362 1409 362 1 outb2
rlabel polycontact 1453 411 1453 411 1 outb2
rlabel ndcontact 1450 396 1450 396 1 s1_bar
rlabel polycontact 1481 404 1481 404 1 s1_bar
rlabel metal1 1492 404 1492 404 7 s1
rlabel ndcontact 1488 396 1488 396 1 s1
rlabel pdcontact 1488 421 1488 421 1 s1
rlabel pdcontact 1460 441 1460 441 1 s1_bar
rlabel pdcontact 1440 441 1440 441 1 vdd
rlabel polycontact 1445 418 1445 418 1 outb1
rlabel ndcontact 1409 440 1409 440 1 outb1
rlabel pdcontact 1409 482 1409 482 1 outb1
rlabel polycontact 1399 467 1399 467 1 b1n
rlabel pdcontact 1365 482 1365 482 1 b1n
rlabel ndcontact 1377 443 1377 443 1 b1n
rlabel ndiffusion 1365 443 1365 443 1 b1m
rlabel polycontact 1368 460 1368 460 1 p1
rlabel polycontact 1356 463 1356 463 1 c1_bar
rlabel ndcontact 1329 439 1329 439 1 c1_bar
rlabel pdcontact 1329 464 1329 464 1 c1_bar
rlabel polycontact 1322 220 1322 220 1 p2
rlabel ndcontact 1329 212 1329 212 1 p2_bar
rlabel pdcontact 1329 237 1329 237 1 p2_bar
rlabel polycontact 1356 216 1356 216 1 p2_bar
rlabel polycontact 1368 209 1368 209 1 c2
rlabel polycontact 1322 280 1322 280 1 c2
rlabel polycontact 1368 293 1368 293 1 p2
rlabel pdcontact 1365 315 1365 315 1 c1n
rlabel ndcontact 1377 276 1377 276 1 c1n
rlabel ndiffusion 1365 276 1365 276 1 c1m
rlabel polycontact 1399 300 1399 300 1 c1n
rlabel pdcontact 1409 315 1409 315 1 outc1
rlabel ndcontact 1409 273 1409 273 1 outc1
rlabel polycontact 1445 251 1445 251 1 outc1
rlabel pdcontact 1440 274 1440 274 1 vdd
rlabel polycontact 1453 244 1453 244 1 outc2
rlabel pdcontact 1460 274 1460 274 1 s2_bar
rlabel polycontact 1481 237 1481 237 1 s2_bar
rlabel ndcontact 1450 229 1450 229 1 s2_bar
rlabel metal1 1492 237 1492 237 7 s2
rlabel pdcontact 1365 237 1365 237 1 c2n
rlabel ndiffusion 1365 198 1365 198 1 c2m
rlabel ndcontact 1377 198 1377 198 1 c2n
rlabel polycontact 1399 220 1399 220 1 c2n
rlabel ndcontact 1409 195 1409 195 1 outc2
rlabel pdcontact 1409 237 1409 237 1 outc2
rlabel polycontact 1323 55 1323 55 1 p3
rlabel ndcontact 1330 47 1330 47 1 p3_bar
rlabel pdcontact 1330 72 1330 72 1 p3_bar
rlabel polycontact 1357 51 1357 51 1 p3_bar
rlabel polycontact 1369 44 1369 44 1 c3
rlabel polycontact 1323 115 1323 115 1 c3
rlabel polycontact 1369 128 1369 128 1 p3
rlabel pdcontact 1366 150 1366 150 1 d1n
rlabel ndcontact 1378 111 1378 111 1 d1n
rlabel ndiffusion 1366 111 1366 111 1 d1m
rlabel polycontact 1400 135 1400 135 1 d1n
rlabel pdcontact 1410 150 1410 150 1 outd1
rlabel ndcontact 1410 108 1410 108 1 outd1
rlabel polycontact 1446 86 1446 86 1 outd1
rlabel polycontact 1454 79 1454 79 1 outd2
rlabel pdcontact 1441 109 1441 109 1 vdd
rlabel pdcontact 1461 109 1461 109 1 s3_bar
rlabel polycontact 1482 72 1482 72 1 s3_bar
rlabel metal1 1493 72 1493 72 7 s3
rlabel pdcontact 1489 89 1489 89 1 s3
rlabel ndcontact 1451 64 1451 64 1 s3_bar
rlabel pdcontact 1366 72 1366 72 1 d2n
rlabel ndcontact 1378 33 1378 33 1 d2n
rlabel ndiffusion 1366 33 1366 33 1 d2m
rlabel polycontact 1400 55 1400 55 1 d2n
rlabel pdcontact 1410 72 1410 72 1 outd2
rlabel ndcontact 1410 30 1410 30 1 outd2
rlabel pdiffusion 1451 110 1451 110 1 dps
rlabel pdiffusion 1450 274 1450 274 1 cps
rlabel pdiffusion 1450 442 1450 442 1 bps
rlabel pdiffusion 1450 604 1450 604 1 aps
rlabel ndcontact 1488 229 1488 229 1 s2
rlabel pdcontact 1488 254 1488 254 1 s2
rlabel ndcontact 1489 64 1489 64 1 s3
rlabel ndcontact 1329 603 1329 603 1 c0_bar
rlabel ndcontact 1329 543 1329 543 1 p0_bar
rlabel pdcontact 1321 568 1321 568 1 vdd
rlabel ndcontact 1321 543 1321 543 1 gnd
rlabel ndcontact 1352 529 1352 529 1 gnd
rlabel pdcontact 1355 568 1355 568 1 vdd
rlabel pdcontact 1375 568 1375 568 1 vdd
rlabel ndcontact 1395 526 1395 526 1 gnd
rlabel pdcontact 1395 568 1395 568 1 vdd
rlabel metal1 1188 286 1188 286 5 VDD
rlabel pdcontact 1179 268 1179 268 1 vdd
rlabel metal1 1189 199 1189 199 1 GND
rlabel ndcontact 1197 208 1197 208 1 gnd
rlabel ndcontact 1179 208 1179 208 1 gnd
rlabel ndcontact 1215 208 1215 208 1 gnd
rlabel ndcontact 1242 230 1242 230 1 gnd
rlabel pdcontact 1242 255 1242 255 1 vdd
rlabel metal1 1092 219 1092 219 5 VDD
rlabel metal1 1079 148 1079 148 2 GND
rlabel ndcontact 1079 161 1079 161 3 gnd
rlabel ndcontact 1133 161 1133 161 1 gnd
rlabel pdcontact 1133 207 1133 207 1 vdd
rlabel pdcontact 1104 207 1104 207 1 vdd
rlabel pdcontact 1082 207 1082 207 1 vdd
rlabel metal1 1092 588 1092 588 5 VDD
rlabel metal1 1079 524 1079 524 2 GND
rlabel metal1 1172 516 1172 516 1 GND
rlabel metal1 1171 588 1171 588 5 VDD
rlabel metal1 1092 501 1092 501 5 VDD
rlabel metal1 1079 430 1079 430 2 GND
rlabel ndcontact 1079 443 1079 443 3 gnd
rlabel ndcontact 1133 443 1133 443 1 gnd
rlabel pdcontact 1133 489 1133 489 1 vdd
rlabel pdcontact 1104 489 1104 489 1 vdd
rlabel pdcontact 1082 489 1082 489 1 vdd
rlabel metal1 1092 406 1092 406 5 VDD
rlabel metal1 1079 342 1079 342 2 GND
rlabel metal1 1188 470 1188 470 5 VDD
rlabel metal1 1189 391 1189 391 1 GND
rlabel ndcontact 1228 421 1228 421 1 gnd
rlabel pdcontact 1228 446 1228 446 1 vdd
rlabel ndcontact 1197 400 1197 400 1 gnd
rlabel ndcontact 1179 400 1179 400 1 gnd
rlabel pdcontact 1179 452 1179 452 1 vdd
rlabel metal1 1092 317 1092 317 5 VDD
rlabel pdcontact 1104 305 1104 305 1 vdd
rlabel pdcontact 1082 305 1082 305 1 vdd
rlabel ndcontact 1079 252 1079 252 3 gnd
rlabel metal1 1079 239 1079 239 2 GND
rlabel pdcontact 1140 305 1140 305 1 vdd
rlabel ndcontact 1140 252 1140 252 1 gnd
rlabel pdcontact 1126 305 1126 305 1 vdd
rlabel metal1 1092 126 1092 126 5 VDD
rlabel metal1 1079 62 1079 62 2 GND
rlabel polycontact 1083 555 1083 555 1 g0
rlabel polycontact 1126 559 1126 559 1 p1g0_bar
rlabel polycontact 1167 547 1167 547 1 p1g0
rlabel polycontact 1175 540 1175 540 1 g1
rlabel polycontact 1203 533 1203 533 1 c2_bar
rlabel metal1 1214 533 1214 533 1 c2
rlabel pdcontact 1082 576 1082 576 1 vdd
rlabel pdcontact 1102 576 1102 576 1 vdd
rlabel pdcontact 1092 576 1092 576 1 p1g0_bar
rlabel ndcontact 1104 537 1104 537 1 p1g0_bar
rlabel ndcontact 1079 537 1079 537 3 gnd
rlabel pdcontact 1122 576 1122 576 1 vdd
rlabel pdcontact 1136 576 1136 576 1 p1g0
rlabel ndcontact 1122 534 1122 534 1 gnd
rlabel ndcontact 1136 534 1136 534 1 p1g0
rlabel pdcontact 1162 570 1162 570 1 vdd
rlabel ndcontact 1162 525 1162 525 1 gnd
rlabel ndcontact 1182 525 1182 525 1 gnd
rlabel ndcontact 1172 525 1172 525 1 c2_bar
rlabel pdcontact 1182 570 1182 570 1 c2_bar
rlabel ndcontact 1202 525 1202 525 1 gnd
rlabel ndcontact 1210 525 1210 525 1 c2
rlabel pdcontact 1210 550 1210 550 1 c2
rlabel pdcontact 1202 550 1202 550 1 vdd
rlabel ndiffusion 1092 537 1092 537 1 n1
rlabel pdiffusion 1172 571 1172 571 1 n2
rlabel polycontact 1107 454 1107 454 1 g0
rlabel ndiffusion 1092 443 1092 443 1 n3
rlabel ndiffusion 1104 443 1104 443 1 n4
rlabel polycontact 1137 472 1137 472 1 p2p1g0_bar
rlabel pdcontact 1114 489 1114 489 1 p2p1g0_bar
rlabel pdcontact 1092 489 1092 489 1 p2p1g0_bar
rlabel pdcontact 1147 489 1147 489 1 p2p1g0
rlabel ndcontact 1147 443 1147 443 1 p2p1g0
rlabel ndcontact 1114 443 1114 443 1 p2p1g0_bar
rlabel polycontact 1184 429 1184 429 1 p2p1g0
rlabel pdcontact 1102 394 1102 394 1 vdd
rlabel pdcontact 1122 394 1122 394 1 vdd
rlabel pdcontact 1082 394 1082 394 1 vdd
rlabel polycontact 1095 366 1095 366 1 g1
rlabel polycontact 1126 377 1126 377 1 p2g1_bar
rlabel pdcontact 1092 394 1092 394 1 p2g1_bar
rlabel ndcontact 1104 355 1104 355 1 p2g1_bar
rlabel ndcontact 1079 355 1079 355 3 gnd
rlabel ndcontact 1122 352 1122 352 1 gnd
rlabel pdcontact 1136 394 1136 394 1 p2g1
rlabel ndcontact 1136 352 1136 352 1 p2g1
rlabel polycontact 1192 422 1192 422 1 p2g1
rlabel polycontact 1200 415 1200 415 1 g2
rlabel ndcontact 1236 421 1236 421 1 c3
rlabel pdcontact 1236 446 1236 446 1 c3
rlabel polycontact 1119 263 1119 263 1 g0
rlabel ndiffusion 1092 355 1092 355 1 n5
rlabel pdiffusion 1189 452 1189 452 1 n6
rlabel pdiffusion 1197 452 1197 452 1 n7
rlabel ndiffusion 1092 252 1092 252 1 n8
rlabel ndiffusion 1104 252 1104 252 1 n9
rlabel ndiffusion 1116 252 1116 252 1 n10
rlabel ndcontact 1126 252 1126 252 1 p3p2p1g0_bar
rlabel pdcontact 1116 305 1116 305 1 p3p2p1g0_bar
rlabel pdcontact 1092 305 1092 305 1 p3p2p1g0_bar
rlabel polycontact 1144 288 1144 288 1 p3p2p1g0_bar
rlabel ndcontact 1154 252 1154 252 1 p3p2p1g0
rlabel pdcontact 1154 305 1154 305 1 p3p2p1g0
rlabel polycontact 1184 245 1184 245 1 p3p2p1g0
rlabel polycontact 1107 172 1107 172 1 g1
rlabel ndiffusion 1092 161 1092 161 1 n11
rlabel ndiffusion 1104 161 1104 161 1 n12
rlabel ndcontact 1114 161 1114 161 1 p3p2g1_bar
rlabel pdcontact 1092 207 1092 207 1 p3p2g1_bar
rlabel pdcontact 1114 207 1114 207 1 p3p2g1_bar
rlabel polycontact 1137 190 1137 190 1 p3p2g1_bar
rlabel ndcontact 1147 161 1147 161 1 p3p2g1
rlabel pdcontact 1147 207 1147 207 1 p3p2g1
rlabel polycontact 1192 238 1192 238 1 p3p2g1
rlabel polycontact 1095 86 1095 86 1 g2
rlabel ndcontact 1079 75 1079 75 3 gnd
rlabel ndcontact 1122 72 1122 72 1 gnd
rlabel ndcontact 1104 75 1104 75 1 p3g2_bar
rlabel pdcontact 1082 114 1082 114 1 vdd
rlabel pdcontact 1092 114 1092 114 1 p3g2_bar
rlabel pdcontact 1102 114 1102 114 1 vdd
rlabel polycontact 1126 97 1126 97 1 p3g2_bar
rlabel pdcontact 1122 114 1122 114 1 vdd
rlabel pdcontact 1136 114 1136 114 1 p3g2
rlabel ndcontact 1136 72 1136 72 1 p3g2
rlabel ndiffusion 1092 75 1092 75 1 n13
rlabel polycontact 1208 224 1208 224 1 p3g2
rlabel pdiffusion 1189 269 1189 269 1 n14
rlabel pdiffusion 1197 269 1197 269 1 n15
rlabel pdiffusion 1205 269 1205 269 1 n16
rlabel ndcontact 1189 208 1189 208 1 cout_bar
rlabel ndcontact 1205 208 1205 208 1 cout_bar
rlabel pdcontact 1215 268 1215 268 1 cout_bar
rlabel polycontact 1243 238 1243 238 1 cout_bar
rlabel metal1 1254 238 1254 238 7 cout
rlabel ndcontact 1250 230 1250 230 1 cout
rlabel pdcontact 1250 255 1250 255 1 cout
rlabel polycontact 1095 548 1095 548 1 p1
rlabel polycontact 1095 461 1095 461 1 p1
rlabel polycontact 1107 270 1107 270 1 p1
rlabel polycontact 1083 468 1083 468 1 p2
rlabel polycontact 1083 373 1083 373 1 p2
rlabel polycontact 1095 277 1095 277 1 p2
rlabel polycontact 1095 179 1095 179 1 p2
rlabel polycontact 1083 284 1083 284 1 p3
rlabel polycontact 1083 186 1083 186 1 p3
rlabel polycontact 1083 93 1083 93 1 p3
rlabel metal1 802 654 802 654 5 VDD
rlabel metal1 805 609 805 609 1 GND
rlabel metal1 802 594 802 594 5 VDD
rlabel metal1 805 549 805 549 1 GND
rlabel metal1 846 595 846 595 5 VDD
rlabel metal1 860 531 860 531 1 GND
rlabel metal1 846 673 846 673 5 VDD
rlabel metal1 860 609 860 609 1 GND
rlabel metal1 930 638 930 638 5 VDD
rlabel metal1 931 566 931 566 1 GND
rlabel ndcontact 802 558 802 558 1 GND
rlabel pdcontact 802 583 802 583 1 VDD
rlabel ndcontact 802 618 802 618 1 GND
rlabel pdcontact 802 643 802 643 1 VDD
rlabel ndcontact 833 544 833 544 1 GND
rlabel ndiffusion 846 544 846 544 1 and2m
rlabel ndcontact 858 544 858 544 1 and2n
rlabel pdcontact 836 583 836 583 1 VDD
rlabel pdcontact 846 583 846 583 1 and2n
rlabel pdcontact 856 583 856 583 1 VDD
rlabel ndcontact 833 622 833 622 1 GND
rlabel ndiffusion 846 622 846 622 1 and1m
rlabel ndcontact 858 622 858 622 1 and1n
rlabel pdcontact 836 661 836 661 1 VDD
rlabel pdcontact 856 661 856 661 1 VDD
rlabel pdcontact 846 661 846 661 1 and1n
rlabel polycontact 880 646 880 646 1 and1n
rlabel pdcontact 876 661 876 661 1 VDD
rlabel pdcontact 890 661 890 661 1 outand1
rlabel ndcontact 890 619 890 619 1 outand1
rlabel ndcontact 876 619 876 619 1 GND
rlabel pdcontact 876 583 876 583 1 VDD
rlabel pdcontact 890 583 890 583 1 outand2
rlabel ndcontact 890 541 890 541 1 outand2
rlabel ndcontact 876 541 876 541 1 GND
rlabel polycontact 880 566 880 566 1 and2n
rlabel polycontact 926 597 926 597 1 outand1
rlabel polycontact 934 590 934 590 1 outand2
rlabel ndcontact 921 575 921 575 1 GND
rlabel ndcontact 941 575 941 575 1 GND
rlabel ndcontact 961 575 961 575 1 GND
rlabel pdcontact 961 600 961 600 1 VDD
rlabel metal1 911 492 911 492 2 GND
rlabel metal1 924 556 924 556 5 VDD
rlabel metal1 802 492 802 492 5 VDD
rlabel metal1 805 447 805 447 1 GND
rlabel metal1 802 432 802 432 5 VDD
rlabel metal1 805 387 805 387 1 GND
rlabel metal1 846 433 846 433 5 VDD
rlabel metal1 860 369 860 369 1 GND
rlabel metal1 846 511 846 511 5 VDD
rlabel metal1 860 447 860 447 1 GND
rlabel ndcontact 802 396 802 396 1 GND
rlabel pdcontact 802 421 802 421 1 VDD
rlabel ndcontact 802 456 802 456 1 GND
rlabel pdcontact 802 481 802 481 1 VDD
rlabel ndcontact 833 382 833 382 1 GND
rlabel pdcontact 836 421 836 421 1 VDD
rlabel pdcontact 856 421 856 421 1 VDD
rlabel ndcontact 833 460 833 460 1 GND
rlabel pdcontact 836 499 836 499 1 VDD
rlabel pdcontact 856 499 856 499 1 VDD
rlabel pdcontact 876 499 876 499 1 VDD
rlabel ndcontact 876 457 876 457 1 GND
rlabel pdcontact 876 421 876 421 1 VDD
rlabel ndcontact 876 379 876 379 1 GND
rlabel metal1 927 476 927 476 5 VDD
rlabel metal1 928 404 928 404 1 GND
rlabel ndcontact 918 413 918 413 1 GND
rlabel ndcontact 938 413 938 413 1 GND
rlabel ndcontact 958 413 958 413 1 GND
rlabel pdcontact 958 438 958 438 1 VDD
rlabel metal1 921 394 921 394 5 VDD
rlabel metal1 908 330 908 330 2 GND
rlabel metal1 802 330 802 330 5 VDD
rlabel metal1 805 285 805 285 1 GND
rlabel metal1 802 270 802 270 5 VDD
rlabel metal1 805 225 805 225 1 GND
rlabel metal1 846 271 846 271 5 VDD
rlabel metal1 860 207 860 207 1 GND
rlabel metal1 846 349 846 349 5 VDD
rlabel metal1 860 285 860 285 1 GND
rlabel metal1 930 314 930 314 5 VDD
rlabel metal1 931 242 931 242 1 GND
rlabel ndcontact 802 234 802 234 1 GND
rlabel pdcontact 802 259 802 259 1 VDD
rlabel ndcontact 802 294 802 294 1 GND
rlabel pdcontact 802 319 802 319 1 VDD
rlabel ndcontact 833 220 833 220 1 GND
rlabel pdcontact 836 259 836 259 1 VDD
rlabel pdcontact 856 259 856 259 1 VDD
rlabel ndcontact 833 298 833 298 1 GND
rlabel pdcontact 836 337 836 337 1 VDD
rlabel pdcontact 856 337 856 337 1 VDD
rlabel pdcontact 876 337 876 337 1 VDD
rlabel ndcontact 876 295 876 295 1 GND
rlabel pdcontact 876 259 876 259 1 VDD
rlabel ndcontact 876 217 876 217 1 GND
rlabel ndcontact 921 251 921 251 1 GND
rlabel ndcontact 941 251 941 251 1 GND
rlabel ndcontact 961 251 961 251 1 GND
rlabel pdcontact 961 276 961 276 1 VDD
rlabel metal1 911 168 911 168 2 GND
rlabel metal1 924 232 924 232 5 VDD
rlabel metal1 802 168 802 168 5 VDD
rlabel metal1 805 123 805 123 1 GND
rlabel metal1 802 108 802 108 5 VDD
rlabel metal1 805 63 805 63 1 GND
rlabel metal1 846 109 846 109 5 VDD
rlabel metal1 860 45 860 45 1 GND
rlabel metal1 846 187 846 187 5 VDD
rlabel metal1 860 123 860 123 1 GND
rlabel ndcontact 802 72 802 72 1 GND
rlabel pdcontact 802 97 802 97 1 VDD
rlabel ndcontact 802 132 802 132 1 GND
rlabel pdcontact 802 157 802 157 1 VDD
rlabel ndcontact 833 58 833 58 1 GND
rlabel pdcontact 836 97 836 97 1 VDD
rlabel pdcontact 856 97 856 97 1 VDD
rlabel ndcontact 833 136 833 136 1 GND
rlabel pdcontact 836 175 836 175 1 VDD
rlabel pdcontact 856 175 856 175 1 VDD
rlabel pdcontact 876 175 876 175 1 VDD
rlabel ndcontact 876 133 876 133 1 GND
rlabel pdcontact 876 97 876 97 1 VDD
rlabel ndcontact 876 55 876 55 1 GND
rlabel metal1 927 152 927 152 5 VDD
rlabel metal1 928 80 928 80 1 GND
rlabel ndcontact 918 89 918 89 1 GND
rlabel ndcontact 938 89 938 89 1 GND
rlabel ndcontact 958 89 958 89 1 GND
rlabel pdcontact 958 114 958 114 1 VDD
rlabel metal1 921 70 921 70 5 VDD
rlabel metal1 908 6 908 6 2 GND
rlabel ndcontact 968 502 968 502 1 g0
rlabel pdcontact 968 544 968 544 1 g0
rlabel ndcontact 954 502 954 502 1 gnd
rlabel ndcontact 936 505 936 505 1 g0_bar
rlabel polycontact 958 527 958 527 1 g0_bar
rlabel pdcontact 924 544 924 544 1 g0_bar
rlabel pdcontact 954 544 954 544 1 vdd
rlabel pdcontact 934 544 934 544 1 vdd
rlabel pdcontact 914 544 914 544 1 vdd
rlabel ndcontact 911 505 911 505 1 gnd
rlabel ndiffusion 923 505 923 505 1 and0m
rlabel polycontact 927 516 927 516 1 b0
rlabel ndcontact 969 575 969 575 1 p0
rlabel metal1 973 583 973 583 7 p0
rlabel pdcontact 969 600 969 600 1 p0
rlabel polycontact 962 583 962 583 1 p0_bar
rlabel ndcontact 931 575 931 575 1 p0_bar
rlabel pdcontact 941 620 941 620 1 p0_bar
rlabel pdcontact 921 620 921 620 1 vdd
rlabel polycontact 803 566 803 566 1 a0
rlabel ndcontact 810 558 810 558 1 a0_bar
rlabel pdcontact 810 583 810 583 1 a0_bar
rlabel polycontact 837 562 837 562 1 a0_bar
rlabel polycontact 849 555 849 555 1 b0
rlabel polycontact 803 626 803 626 1 b0
rlabel pdcontact 810 643 810 643 1 b0_bar
rlabel ndcontact 810 618 810 618 1 b0_bar
rlabel polycontact 837 642 837 642 1 b0_bar
rlabel polycontact 849 639 849 639 1 a0
rlabel polycontact 915 523 915 523 1 a0
rlabel ndcontact 951 340 951 340 1 gnd
rlabel ndcontact 965 340 965 340 1 g1
rlabel pdcontact 965 382 965 382 1 g1
rlabel pdcontact 951 382 951 382 1 vdd
rlabel polycontact 955 365 955 365 1 g1_bar
rlabel ndcontact 933 343 933 343 1 g1_bar
rlabel ndcontact 908 343 908 343 1 gnd
rlabel pdcontact 921 382 921 382 1 g1_bar
rlabel pdcontact 931 382 931 382 1 vdd
rlabel pdcontact 911 382 911 382 1 vdd
rlabel polycontact 924 354 924 354 1 b1
rlabel polycontact 912 361 912 361 1 a1
rlabel ndcontact 966 413 966 413 1 p1
rlabel pdcontact 966 438 966 438 1 p1
rlabel polycontact 959 421 959 421 1 p1_bar
rlabel ndcontact 928 413 928 413 1 p1_bar
rlabel pdcontact 938 458 938 458 1 p1_bar
rlabel pdcontact 918 458 918 458 1 vdd
rlabel polycontact 803 404 803 404 1 a1
rlabel ndcontact 810 396 810 396 1 a1_bar
rlabel pdcontact 810 421 810 421 1 a1_bar
rlabel polycontact 837 400 837 400 1 a1_bar
rlabel polycontact 849 393 849 393 1 b1
rlabel polycontact 803 464 803 464 1 b1
rlabel ndcontact 810 456 810 456 1 b1_bar
rlabel pdcontact 810 481 810 481 1 b1_bar
rlabel polycontact 837 480 837 480 1 b1_bar
rlabel polycontact 849 477 849 477 1 a1
rlabel metal1 972 203 972 203 7 g2
rlabel ndcontact 968 178 968 178 1 g2
rlabel pdcontact 968 220 968 220 1 g2
rlabel ndcontact 954 178 954 178 1 gnd
rlabel ndcontact 936 181 936 181 1 g2_bar
rlabel ndcontact 911 181 911 181 1 gnd
rlabel polycontact 958 203 958 203 1 g2_bar
rlabel polycontact 927 192 927 192 1 b2
rlabel polycontact 915 199 915 199 1 a2
rlabel pdcontact 954 220 954 220 1 vdd
rlabel pdcontact 934 220 934 220 1 vdd
rlabel pdcontact 914 220 914 220 1 vdd
rlabel pdcontact 924 220 924 220 1 g2_bar
rlabel polycontact 962 259 962 259 1 p2_bar
rlabel ndcontact 931 251 931 251 1 p2_bar
rlabel pdcontact 941 295 941 295 1 p2_bar
rlabel pdcontact 921 296 921 296 1 vdd
rlabel polycontact 803 242 803 242 1 a2
rlabel ndcontact 810 234 810 234 1 a2_bar
rlabel pdcontact 810 259 810 259 1 a2_bar
rlabel polycontact 837 238 837 238 1 a2_bar
rlabel polycontact 849 231 849 231 1 b2
rlabel polycontact 803 302 803 302 1 b2
rlabel pdcontact 810 319 810 319 1 b2_bar
rlabel ndcontact 810 294 810 294 1 b2_bar
rlabel polycontact 837 318 837 318 1 b2_bar
rlabel polycontact 849 315 849 315 1 a2
rlabel ndcontact 951 16 951 16 1 gnd
rlabel ndcontact 965 16 965 16 1 g3
rlabel pdcontact 965 58 965 58 1 g3
rlabel pdcontact 951 58 951 58 1 vdd
rlabel polycontact 955 41 955 41 1 g3_bar
rlabel ndcontact 933 19 933 19 1 g3_bar
rlabel ndcontact 908 19 908 19 1 gnd
rlabel polycontact 924 30 924 30 1 b3
rlabel polycontact 912 37 912 37 1 a3
rlabel pdcontact 931 58 931 58 1 vdd
rlabel pdcontact 911 58 911 58 1 vdd
rlabel pdcontact 921 58 921 58 1 g3_bar
rlabel ndcontact 966 89 966 89 1 p3
rlabel metal1 970 97 970 97 1 p3
rlabel pdcontact 966 114 966 114 1 p3
rlabel polycontact 959 97 959 97 1 p3_bar
rlabel ndcontact 928 89 928 89 1 p3_bar
rlabel pdcontact 938 134 938 134 1 p3_bar
rlabel pdcontact 918 134 918 134 1 vdd
rlabel polycontact 803 80 803 80 1 a3
rlabel ndcontact 810 72 810 72 1 a3_bar
rlabel pdcontact 810 97 810 97 1 a3_bar
rlabel polycontact 837 76 837 76 1 a3_bar
rlabel polycontact 849 69 849 69 1 b3
rlabel polycontact 803 140 803 140 1 b3
rlabel pdcontact 810 157 810 157 1 b3_bar
rlabel ndcontact 810 132 810 132 1 b3_bar
rlabel polycontact 837 156 837 156 1 b3_bar
rlabel polycontact 849 153 849 153 1 a3
rlabel polycontact 1200 231 1200 231 1 g3
rlabel pdcontact 969 276 969 276 1 p2
rlabel ndcontact 969 251 969 251 1 p2
rlabel ndiffusion 846 460 846 460 1 anda1m
rlabel ndcontact 858 460 858 460 1 anda1n
rlabel pdcontact 846 499 846 499 1 anda1n
rlabel polycontact 880 484 880 484 1 anda1n
rlabel pdcontact 890 499 890 499 1 outanda1
rlabel ndcontact 890 457 890 457 1 outanda1
rlabel polycontact 923 435 923 435 1 outanda1
rlabel pdcontact 846 421 846 421 1 anda2n
rlabel ndcontact 858 382 858 382 1 anda2n
rlabel ndiffusion 846 382 846 382 1 anda2m
rlabel polycontact 880 404 880 404 1 anda2n
rlabel pdcontact 890 421 890 421 1 outanda2
rlabel ndcontact 890 379 890 379 1 outanda2
rlabel polycontact 931 428 931 428 1 outanda2
rlabel pdcontact 846 337 846 337 1 andb1n
rlabel ndiffusion 846 298 846 298 1 andb1m
rlabel ndcontact 858 298 858 298 1 andb1n
rlabel polycontact 880 322 880 322 1 andb1n
rlabel pdcontact 890 337 890 337 1 outband1
rlabel ndcontact 890 295 890 295 1 outband1
rlabel polycontact 926 273 926 273 1 outband1
rlabel pdcontact 846 259 846 259 1 andb2n
rlabel polycontact 880 242 880 242 1 andb2n
rlabel ndcontact 858 220 858 220 1 andb2n
rlabel ndiffusion 846 220 846 220 1 andb2m
rlabel pdcontact 890 259 890 259 1 outband2
rlabel ndcontact 890 217 890 217 1 outband2
rlabel polycontact 934 266 934 266 1 outband2
rlabel pdcontact 846 175 846 175 1 andc1n
rlabel polycontact 880 160 880 160 1 andc1n
rlabel ndcontact 858 136 858 136 1 andc1n
rlabel ndiffusion 846 136 846 136 1 andc1m
rlabel pdcontact 890 175 890 175 1 outcand1
rlabel ndcontact 890 133 890 133 1 outcand1
rlabel polycontact 923 111 923 111 1 outcand1
rlabel pdcontact 846 97 846 97 1 andc2n
rlabel ndcontact 858 58 858 58 1 andc2n
rlabel polycontact 880 80 880 80 1 andc2n
rlabel ndiffusion 846 58 846 58 1 andc2m
rlabel ndcontact 890 55 890 55 1 outcand2
rlabel pdcontact 890 97 890 97 1 outcand2
rlabel polycontact 931 104 931 104 1 outcand2
rlabel polycontact 1368 376 1368 376 1 g0
rlabel polycontact 1322 447 1322 447 1 g0
rlabel pdcontact 1207 452 1207 452 1 c3_bar
rlabel ndcontact 1207 400 1207 400 1 c3_bar
rlabel ndcontact 1189 400 1189 400 1 c3_bar
rlabel polycontact 1229 429 1229 429 1 c3_bar
rlabel ndcontact 1330 107 1330 107 1 c3_bar1
rlabel pdcontact 1330 132 1330 132 1 c3_bar1
rlabel polycontact 1357 131 1357 131 1 c3_bar1
rlabel polycontact 1356 296 1356 296 1 c2_bar1
rlabel ndcontact 1329 272 1329 272 1 c2_bar1
rlabel pdcontact 1329 297 1329 297 1 c2_bar1
<< end >>
