magic
tech scmos
timestamp 1732013933
<< nwell >>
rect 18 102 42 126
rect 52 120 122 144
rect 137 85 173 109
rect 137 73 201 85
rect 18 42 42 66
rect 52 42 122 66
rect 177 59 201 73
rect 18 -62 42 -38
rect 52 -44 122 -20
rect 137 -79 173 -55
rect 137 -91 201 -79
rect 18 -122 42 -98
rect 52 -122 122 -98
rect 177 -105 201 -91
rect 18 -229 42 -205
rect 52 -211 122 -187
rect 137 -246 173 -222
rect 137 -258 201 -246
rect 18 -289 42 -265
rect 52 -289 122 -265
rect 177 -272 201 -258
rect 19 -394 43 -370
rect 53 -376 123 -352
rect 138 -411 174 -387
rect 138 -423 202 -411
rect 19 -454 43 -430
rect 53 -454 123 -430
rect 178 -437 202 -423
<< ntransistor >>
rect 29 86 31 92
rect 63 87 65 99
rect 75 87 77 99
rect 106 87 108 93
rect 29 26 31 32
rect 63 9 65 21
rect 75 9 77 21
rect 150 43 152 49
rect 158 43 160 49
rect 188 43 190 49
rect 106 9 108 15
rect 29 -78 31 -72
rect 63 -77 65 -65
rect 75 -77 77 -65
rect 106 -77 108 -71
rect 29 -138 31 -132
rect 63 -155 65 -143
rect 75 -155 77 -143
rect 150 -121 152 -115
rect 158 -121 160 -115
rect 188 -121 190 -115
rect 106 -155 108 -149
rect 29 -245 31 -239
rect 63 -244 65 -232
rect 75 -244 77 -232
rect 106 -244 108 -238
rect 29 -305 31 -299
rect 63 -322 65 -310
rect 75 -322 77 -310
rect 150 -288 152 -282
rect 158 -288 160 -282
rect 188 -288 190 -282
rect 106 -322 108 -316
rect 30 -410 32 -404
rect 64 -409 66 -397
rect 76 -409 78 -397
rect 107 -409 109 -403
rect 30 -470 32 -464
rect 64 -487 66 -475
rect 76 -487 78 -475
rect 151 -453 153 -447
rect 159 -453 161 -447
rect 189 -453 191 -447
rect 107 -487 109 -481
<< ptransistor >>
rect 63 126 65 138
rect 75 126 77 138
rect 106 126 108 138
rect 29 108 31 120
rect 150 79 152 103
rect 158 79 160 103
rect 29 48 31 60
rect 63 48 65 60
rect 75 48 77 60
rect 106 48 108 60
rect 188 65 190 77
rect 63 -38 65 -26
rect 75 -38 77 -26
rect 106 -38 108 -26
rect 29 -56 31 -44
rect 150 -85 152 -61
rect 158 -85 160 -61
rect 29 -116 31 -104
rect 63 -116 65 -104
rect 75 -116 77 -104
rect 106 -116 108 -104
rect 188 -99 190 -87
rect 63 -205 65 -193
rect 75 -205 77 -193
rect 106 -205 108 -193
rect 29 -223 31 -211
rect 150 -252 152 -228
rect 158 -252 160 -228
rect 29 -283 31 -271
rect 63 -283 65 -271
rect 75 -283 77 -271
rect 106 -283 108 -271
rect 188 -266 190 -254
rect 64 -370 66 -358
rect 76 -370 78 -358
rect 107 -370 109 -358
rect 30 -388 32 -376
rect 151 -417 153 -393
rect 159 -417 161 -393
rect 30 -448 32 -436
rect 64 -448 66 -436
rect 76 -448 78 -436
rect 107 -448 109 -436
rect 189 -431 191 -419
<< ndiffusion >>
rect 28 86 29 92
rect 31 86 32 92
rect 59 87 63 99
rect 65 87 75 99
rect 77 87 80 99
rect 102 87 106 93
rect 108 87 112 93
rect 28 26 29 32
rect 31 26 32 32
rect 59 9 63 21
rect 65 9 75 21
rect 77 9 80 21
rect 147 43 150 49
rect 152 43 153 49
rect 157 43 158 49
rect 160 43 163 49
rect 187 43 188 49
rect 190 43 191 49
rect 102 9 106 15
rect 108 9 112 15
rect 28 -78 29 -72
rect 31 -78 32 -72
rect 59 -77 63 -65
rect 65 -77 75 -65
rect 77 -77 80 -65
rect 102 -77 106 -71
rect 108 -77 112 -71
rect 28 -138 29 -132
rect 31 -138 32 -132
rect 59 -155 63 -143
rect 65 -155 75 -143
rect 77 -155 80 -143
rect 147 -121 150 -115
rect 152 -121 153 -115
rect 157 -121 158 -115
rect 160 -121 163 -115
rect 187 -121 188 -115
rect 190 -121 191 -115
rect 102 -155 106 -149
rect 108 -155 112 -149
rect 28 -245 29 -239
rect 31 -245 32 -239
rect 59 -244 63 -232
rect 65 -244 75 -232
rect 77 -244 80 -232
rect 102 -244 106 -238
rect 108 -244 112 -238
rect 28 -305 29 -299
rect 31 -305 32 -299
rect 59 -322 63 -310
rect 65 -322 75 -310
rect 77 -322 80 -310
rect 147 -288 150 -282
rect 152 -288 153 -282
rect 157 -288 158 -282
rect 160 -288 163 -282
rect 187 -288 188 -282
rect 190 -288 191 -282
rect 102 -322 106 -316
rect 108 -322 112 -316
rect 29 -410 30 -404
rect 32 -410 33 -404
rect 60 -409 64 -397
rect 66 -409 76 -397
rect 78 -409 81 -397
rect 103 -409 107 -403
rect 109 -409 113 -403
rect 29 -470 30 -464
rect 32 -470 33 -464
rect 60 -487 64 -475
rect 66 -487 76 -475
rect 78 -487 81 -475
rect 148 -453 151 -447
rect 153 -453 154 -447
rect 158 -453 159 -447
rect 161 -453 164 -447
rect 188 -453 189 -447
rect 191 -453 192 -447
rect 103 -487 107 -481
rect 109 -487 113 -481
<< pdiffusion >>
rect 62 126 63 138
rect 65 126 68 138
rect 72 126 75 138
rect 77 126 78 138
rect 102 126 106 138
rect 108 126 112 138
rect 28 108 29 120
rect 31 108 32 120
rect 147 79 150 103
rect 152 79 158 103
rect 160 79 163 103
rect 28 48 29 60
rect 31 48 32 60
rect 62 48 63 60
rect 65 48 68 60
rect 72 48 75 60
rect 77 48 78 60
rect 102 48 106 60
rect 108 48 112 60
rect 187 65 188 77
rect 190 65 191 77
rect 62 -38 63 -26
rect 65 -38 68 -26
rect 72 -38 75 -26
rect 77 -38 78 -26
rect 102 -38 106 -26
rect 108 -38 112 -26
rect 28 -56 29 -44
rect 31 -56 32 -44
rect 147 -85 150 -61
rect 152 -85 158 -61
rect 160 -85 163 -61
rect 28 -116 29 -104
rect 31 -116 32 -104
rect 62 -116 63 -104
rect 65 -116 68 -104
rect 72 -116 75 -104
rect 77 -116 78 -104
rect 102 -116 106 -104
rect 108 -116 112 -104
rect 187 -99 188 -87
rect 190 -99 191 -87
rect 62 -205 63 -193
rect 65 -205 68 -193
rect 72 -205 75 -193
rect 77 -205 78 -193
rect 102 -205 106 -193
rect 108 -205 112 -193
rect 28 -223 29 -211
rect 31 -223 32 -211
rect 147 -252 150 -228
rect 152 -252 158 -228
rect 160 -252 163 -228
rect 28 -283 29 -271
rect 31 -283 32 -271
rect 62 -283 63 -271
rect 65 -283 68 -271
rect 72 -283 75 -271
rect 77 -283 78 -271
rect 102 -283 106 -271
rect 108 -283 112 -271
rect 187 -266 188 -254
rect 190 -266 191 -254
rect 63 -370 64 -358
rect 66 -370 69 -358
rect 73 -370 76 -358
rect 78 -370 79 -358
rect 103 -370 107 -358
rect 109 -370 113 -358
rect 29 -388 30 -376
rect 32 -388 33 -376
rect 148 -417 151 -393
rect 153 -417 159 -393
rect 161 -417 164 -393
rect 29 -448 30 -436
rect 32 -448 33 -436
rect 63 -448 64 -436
rect 66 -448 69 -436
rect 73 -448 76 -436
rect 78 -448 79 -436
rect 103 -448 107 -436
rect 109 -448 113 -436
rect 188 -431 189 -419
rect 191 -431 192 -419
<< ndcontact >>
rect 24 86 28 92
rect 32 86 36 92
rect 55 87 59 99
rect 80 87 84 99
rect 98 87 102 93
rect 112 87 116 93
rect 24 26 28 32
rect 32 26 36 32
rect 55 9 59 21
rect 80 9 84 21
rect 143 43 147 49
rect 153 43 157 49
rect 163 43 167 49
rect 183 43 187 49
rect 191 43 195 49
rect 98 9 102 15
rect 112 9 116 15
rect 24 -78 28 -72
rect 32 -78 36 -72
rect 55 -77 59 -65
rect 80 -77 84 -65
rect 98 -77 102 -71
rect 112 -77 116 -71
rect 24 -138 28 -132
rect 32 -138 36 -132
rect 55 -155 59 -143
rect 80 -155 84 -143
rect 143 -121 147 -115
rect 153 -121 157 -115
rect 163 -121 167 -115
rect 183 -121 187 -115
rect 191 -121 195 -115
rect 98 -155 102 -149
rect 112 -155 116 -149
rect 24 -245 28 -239
rect 32 -245 36 -239
rect 55 -244 59 -232
rect 80 -244 84 -232
rect 98 -244 102 -238
rect 112 -244 116 -238
rect 24 -305 28 -299
rect 32 -305 36 -299
rect 55 -322 59 -310
rect 80 -322 84 -310
rect 143 -288 147 -282
rect 153 -288 157 -282
rect 163 -288 167 -282
rect 183 -288 187 -282
rect 191 -288 195 -282
rect 98 -322 102 -316
rect 112 -322 116 -316
rect 25 -410 29 -404
rect 33 -410 37 -404
rect 56 -409 60 -397
rect 81 -409 85 -397
rect 99 -409 103 -403
rect 113 -409 117 -403
rect 25 -470 29 -464
rect 33 -470 37 -464
rect 56 -487 60 -475
rect 81 -487 85 -475
rect 144 -453 148 -447
rect 154 -453 158 -447
rect 164 -453 168 -447
rect 184 -453 188 -447
rect 192 -453 196 -447
rect 99 -487 103 -481
rect 113 -487 117 -481
<< pdcontact >>
rect 58 126 62 138
rect 68 126 72 138
rect 78 126 82 138
rect 98 126 102 138
rect 112 126 116 138
rect 24 108 28 120
rect 32 108 36 120
rect 143 79 147 103
rect 163 79 167 103
rect 24 48 28 60
rect 32 48 36 60
rect 58 48 62 60
rect 68 48 72 60
rect 78 48 82 60
rect 98 48 102 60
rect 112 48 116 60
rect 183 65 187 77
rect 191 65 195 77
rect 58 -38 62 -26
rect 68 -38 72 -26
rect 78 -38 82 -26
rect 98 -38 102 -26
rect 112 -38 116 -26
rect 24 -56 28 -44
rect 32 -56 36 -44
rect 143 -85 147 -61
rect 163 -85 167 -61
rect 24 -116 28 -104
rect 32 -116 36 -104
rect 58 -116 62 -104
rect 68 -116 72 -104
rect 78 -116 82 -104
rect 98 -116 102 -104
rect 112 -116 116 -104
rect 183 -99 187 -87
rect 191 -99 195 -87
rect 58 -205 62 -193
rect 68 -205 72 -193
rect 78 -205 82 -193
rect 98 -205 102 -193
rect 112 -205 116 -193
rect 24 -223 28 -211
rect 32 -223 36 -211
rect 143 -252 147 -228
rect 163 -252 167 -228
rect 24 -283 28 -271
rect 32 -283 36 -271
rect 58 -283 62 -271
rect 68 -283 72 -271
rect 78 -283 82 -271
rect 98 -283 102 -271
rect 112 -283 116 -271
rect 183 -266 187 -254
rect 191 -266 195 -254
rect 59 -370 63 -358
rect 69 -370 73 -358
rect 79 -370 83 -358
rect 99 -370 103 -358
rect 113 -370 117 -358
rect 25 -388 29 -376
rect 33 -388 37 -376
rect 144 -417 148 -393
rect 164 -417 168 -393
rect 25 -448 29 -436
rect 33 -448 37 -436
rect 59 -448 63 -436
rect 69 -448 73 -436
rect 79 -448 83 -436
rect 99 -448 103 -436
rect 113 -448 117 -436
rect 184 -431 188 -419
rect 192 -431 196 -419
<< polysilicon >>
rect 63 138 65 141
rect 75 138 77 141
rect 106 138 108 141
rect 29 120 31 123
rect 29 92 31 108
rect 63 99 65 126
rect 75 99 77 126
rect 106 93 108 126
rect 150 103 152 106
rect 158 103 160 106
rect 29 83 31 86
rect 63 84 65 87
rect 75 84 77 87
rect 106 84 108 87
rect 150 70 152 79
rect 29 60 31 63
rect 63 60 65 63
rect 75 60 77 63
rect 106 60 108 63
rect 150 49 152 66
rect 158 63 160 79
rect 188 77 190 80
rect 158 49 160 59
rect 188 49 190 65
rect 29 32 31 48
rect 29 23 31 26
rect 63 21 65 48
rect 75 21 77 48
rect 106 15 108 48
rect 150 40 152 43
rect 158 40 160 43
rect 188 39 190 43
rect 63 6 65 9
rect 75 6 77 9
rect 106 6 108 9
rect 63 -26 65 -23
rect 75 -26 77 -23
rect 106 -26 108 -23
rect 29 -44 31 -41
rect 29 -72 31 -56
rect 63 -65 65 -38
rect 75 -65 77 -38
rect 106 -71 108 -38
rect 150 -61 152 -58
rect 158 -61 160 -58
rect 29 -81 31 -78
rect 63 -80 65 -77
rect 75 -80 77 -77
rect 106 -80 108 -77
rect 150 -94 152 -85
rect 29 -104 31 -101
rect 63 -104 65 -101
rect 75 -104 77 -101
rect 106 -104 108 -101
rect 150 -115 152 -98
rect 158 -101 160 -85
rect 188 -87 190 -84
rect 158 -115 160 -105
rect 188 -115 190 -99
rect 29 -132 31 -116
rect 29 -141 31 -138
rect 63 -143 65 -116
rect 75 -143 77 -116
rect 106 -149 108 -116
rect 150 -124 152 -121
rect 158 -124 160 -121
rect 188 -125 190 -121
rect 63 -158 65 -155
rect 75 -158 77 -155
rect 106 -158 108 -155
rect 63 -193 65 -190
rect 75 -193 77 -190
rect 106 -193 108 -190
rect 29 -211 31 -208
rect 29 -239 31 -223
rect 63 -232 65 -205
rect 75 -232 77 -205
rect 106 -238 108 -205
rect 150 -228 152 -225
rect 158 -228 160 -225
rect 29 -248 31 -245
rect 63 -247 65 -244
rect 75 -247 77 -244
rect 106 -247 108 -244
rect 150 -261 152 -252
rect 29 -271 31 -268
rect 63 -271 65 -268
rect 75 -271 77 -268
rect 106 -271 108 -268
rect 150 -282 152 -265
rect 158 -268 160 -252
rect 188 -254 190 -251
rect 158 -282 160 -272
rect 188 -282 190 -266
rect 29 -299 31 -283
rect 29 -308 31 -305
rect 63 -310 65 -283
rect 75 -310 77 -283
rect 106 -316 108 -283
rect 150 -291 152 -288
rect 158 -291 160 -288
rect 188 -292 190 -288
rect 63 -325 65 -322
rect 75 -325 77 -322
rect 106 -325 108 -322
rect 64 -358 66 -355
rect 76 -358 78 -355
rect 107 -358 109 -355
rect 30 -376 32 -373
rect 30 -404 32 -388
rect 64 -397 66 -370
rect 76 -397 78 -370
rect 107 -403 109 -370
rect 151 -393 153 -390
rect 159 -393 161 -390
rect 30 -413 32 -410
rect 64 -412 66 -409
rect 76 -412 78 -409
rect 107 -412 109 -409
rect 151 -426 153 -417
rect 30 -436 32 -433
rect 64 -436 66 -433
rect 76 -436 78 -433
rect 107 -436 109 -433
rect 151 -447 153 -430
rect 159 -433 161 -417
rect 189 -419 191 -416
rect 159 -447 161 -437
rect 189 -447 191 -431
rect 30 -464 32 -448
rect 30 -473 32 -470
rect 64 -475 66 -448
rect 76 -475 78 -448
rect 107 -481 109 -448
rect 151 -456 153 -453
rect 159 -456 161 -453
rect 189 -457 191 -453
rect 64 -490 66 -487
rect 76 -490 78 -487
rect 107 -490 109 -487
<< polycontact >>
rect 59 111 63 115
rect 25 95 29 99
rect 71 108 75 112
rect 102 115 106 119
rect 148 66 152 70
rect 156 59 160 63
rect 184 52 188 56
rect 25 35 29 39
rect 59 31 63 35
rect 71 24 75 28
rect 102 35 106 39
rect 59 -53 63 -49
rect 25 -69 29 -65
rect 71 -56 75 -52
rect 102 -49 106 -45
rect 148 -98 152 -94
rect 156 -105 160 -101
rect 184 -112 188 -108
rect 25 -129 29 -125
rect 59 -133 63 -129
rect 71 -140 75 -136
rect 102 -129 106 -125
rect 59 -220 63 -216
rect 25 -236 29 -232
rect 71 -223 75 -219
rect 102 -216 106 -212
rect 148 -265 152 -261
rect 156 -272 160 -268
rect 184 -279 188 -275
rect 25 -296 29 -292
rect 59 -300 63 -296
rect 71 -307 75 -303
rect 102 -296 106 -292
rect 60 -385 64 -381
rect 26 -401 30 -397
rect 72 -388 76 -384
rect 103 -381 107 -377
rect 149 -430 153 -426
rect 157 -437 161 -433
rect 185 -444 189 -440
rect 26 -461 30 -457
rect 60 -465 64 -461
rect 72 -472 76 -468
rect 103 -461 107 -457
<< metal1 >>
rect 52 142 102 146
rect 58 138 62 142
rect 78 138 82 142
rect 18 124 42 128
rect 98 138 102 142
rect 24 120 28 124
rect 68 119 72 126
rect 68 115 102 119
rect 112 117 116 126
rect 32 99 36 108
rect 46 111 59 115
rect 46 99 50 111
rect 67 106 71 112
rect 60 102 71 106
rect 80 99 84 115
rect 5 95 25 99
rect 32 95 50 99
rect 32 92 36 95
rect 112 113 134 117
rect 112 93 116 113
rect 24 82 28 86
rect 55 82 59 87
rect 98 82 102 87
rect 18 78 42 82
rect 52 78 102 82
rect 130 70 134 113
rect 137 107 176 111
rect 143 103 147 107
rect 172 85 176 107
rect 172 81 187 85
rect 18 64 42 68
rect 52 64 102 68
rect 130 66 148 70
rect 24 60 28 64
rect 58 60 62 64
rect 78 60 82 64
rect 98 60 102 64
rect 32 39 36 48
rect 68 39 72 48
rect 112 39 116 48
rect 130 59 156 63
rect 130 39 134 59
rect 163 56 167 79
rect 183 77 187 81
rect 191 56 195 65
rect 153 52 184 56
rect 191 52 199 56
rect 153 49 157 52
rect 191 49 195 52
rect 143 39 147 43
rect 163 39 167 43
rect 183 39 187 43
rect 14 35 25 39
rect 32 35 54 39
rect 68 35 102 39
rect 112 35 134 39
rect 137 35 187 39
rect 32 32 36 35
rect 50 31 59 35
rect 24 22 28 26
rect 47 24 71 28
rect 18 18 42 22
rect 47 7 51 24
rect 80 21 84 35
rect 112 15 116 35
rect 55 4 59 9
rect 98 4 102 9
rect 52 0 102 4
rect 52 -22 102 -18
rect 58 -26 62 -22
rect 78 -26 82 -22
rect 18 -40 42 -36
rect 98 -26 102 -22
rect 24 -44 28 -40
rect 68 -45 72 -38
rect 68 -49 102 -45
rect 112 -47 116 -38
rect 32 -65 36 -56
rect 46 -53 59 -49
rect 46 -65 50 -53
rect 67 -58 71 -52
rect 60 -62 71 -58
rect 80 -65 84 -49
rect 5 -69 25 -65
rect 32 -69 50 -65
rect 32 -72 36 -69
rect 112 -51 134 -47
rect 112 -71 116 -51
rect 24 -82 28 -78
rect 55 -82 59 -77
rect 98 -82 102 -77
rect 18 -86 42 -82
rect 52 -86 102 -82
rect 130 -94 134 -51
rect 137 -57 176 -53
rect 143 -61 147 -57
rect 172 -79 176 -57
rect 172 -83 187 -79
rect 18 -100 42 -96
rect 52 -100 102 -96
rect 130 -98 148 -94
rect 24 -104 28 -100
rect 58 -104 62 -100
rect 78 -104 82 -100
rect 98 -104 102 -100
rect 32 -125 36 -116
rect 68 -125 72 -116
rect 112 -125 116 -116
rect 130 -105 156 -101
rect 130 -125 134 -105
rect 163 -108 167 -85
rect 183 -87 187 -83
rect 191 -108 195 -99
rect 153 -112 184 -108
rect 191 -112 199 -108
rect 153 -115 157 -112
rect 191 -115 195 -112
rect 143 -125 147 -121
rect 163 -125 167 -121
rect 183 -125 187 -121
rect 14 -129 25 -125
rect 32 -129 54 -125
rect 68 -129 102 -125
rect 112 -129 134 -125
rect 137 -129 187 -125
rect 32 -132 36 -129
rect 50 -133 59 -129
rect 24 -142 28 -138
rect 47 -140 71 -136
rect 18 -146 42 -142
rect 47 -157 51 -140
rect 80 -143 84 -129
rect 112 -149 116 -129
rect 55 -160 59 -155
rect 98 -160 102 -155
rect 52 -163 102 -160
rect 52 -189 102 -185
rect 58 -193 62 -189
rect 78 -193 82 -189
rect 18 -207 42 -203
rect 98 -193 102 -189
rect 24 -211 28 -207
rect 68 -212 72 -205
rect 68 -216 102 -212
rect 112 -214 116 -205
rect 32 -232 36 -223
rect 46 -220 59 -216
rect 46 -232 50 -220
rect 67 -225 71 -219
rect 60 -229 71 -225
rect 80 -232 84 -216
rect 5 -236 25 -232
rect 32 -236 50 -232
rect 32 -239 36 -236
rect 112 -218 134 -214
rect 112 -238 116 -218
rect 24 -249 28 -245
rect 55 -249 59 -244
rect 98 -249 102 -244
rect 18 -253 42 -249
rect 52 -253 102 -249
rect 130 -261 134 -218
rect 137 -224 176 -220
rect 143 -228 147 -224
rect 172 -246 176 -224
rect 172 -250 187 -246
rect 18 -267 42 -263
rect 52 -267 102 -263
rect 130 -265 148 -261
rect 24 -271 28 -267
rect 58 -271 62 -267
rect 78 -271 82 -267
rect 98 -271 102 -267
rect 32 -292 36 -283
rect 68 -292 72 -283
rect 112 -292 116 -283
rect 130 -272 156 -268
rect 130 -292 134 -272
rect 163 -275 167 -252
rect 183 -254 187 -250
rect 191 -275 195 -266
rect 153 -279 184 -275
rect 191 -279 199 -275
rect 153 -282 157 -279
rect 191 -282 195 -279
rect 143 -292 147 -288
rect 163 -292 167 -288
rect 183 -292 187 -288
rect 14 -296 25 -292
rect 32 -296 54 -292
rect 68 -296 102 -292
rect 112 -296 134 -292
rect 137 -296 187 -292
rect 32 -299 36 -296
rect 50 -300 59 -296
rect 24 -309 28 -305
rect 47 -307 71 -303
rect 18 -313 42 -309
rect 47 -324 51 -307
rect 80 -310 84 -296
rect 112 -316 116 -296
rect 55 -327 59 -322
rect 98 -327 102 -322
rect 52 -330 102 -327
rect 53 -354 103 -350
rect 59 -358 63 -354
rect 79 -358 83 -354
rect 19 -372 43 -368
rect 99 -358 103 -354
rect 25 -376 29 -372
rect 69 -377 73 -370
rect 69 -381 103 -377
rect 113 -379 117 -370
rect 33 -397 37 -388
rect 47 -385 60 -381
rect 47 -397 51 -385
rect 68 -390 72 -384
rect 61 -394 72 -390
rect 81 -397 85 -381
rect 6 -401 26 -397
rect 33 -401 51 -397
rect 33 -404 37 -401
rect 113 -383 135 -379
rect 113 -403 117 -383
rect 25 -414 29 -410
rect 56 -414 60 -409
rect 99 -414 103 -409
rect 19 -418 43 -414
rect 53 -418 103 -414
rect 131 -426 135 -383
rect 138 -389 177 -385
rect 144 -393 148 -389
rect 173 -411 177 -389
rect 173 -415 188 -411
rect 19 -432 43 -428
rect 53 -432 103 -428
rect 131 -430 149 -426
rect 25 -436 29 -432
rect 59 -436 63 -432
rect 79 -436 83 -432
rect 99 -436 103 -432
rect 33 -457 37 -448
rect 69 -457 73 -448
rect 113 -457 117 -448
rect 131 -437 157 -433
rect 131 -457 135 -437
rect 164 -440 168 -417
rect 184 -419 188 -415
rect 192 -440 196 -431
rect 154 -444 185 -440
rect 192 -444 200 -440
rect 154 -447 158 -444
rect 192 -447 196 -444
rect 144 -457 148 -453
rect 164 -457 168 -453
rect 184 -457 188 -453
rect 15 -461 26 -457
rect 33 -461 55 -457
rect 69 -461 103 -457
rect 113 -461 135 -457
rect 138 -461 188 -457
rect 33 -464 37 -461
rect 51 -465 60 -461
rect 25 -474 29 -470
rect 48 -472 72 -468
rect 19 -478 43 -474
rect 48 -489 52 -472
rect 81 -475 85 -461
rect 113 -481 117 -461
rect 56 -492 60 -487
rect 99 -492 103 -487
rect 53 -496 103 -492
<< m2contact >>
rect 55 102 60 107
rect 0 94 5 99
rect 9 34 14 39
rect 42 7 47 12
rect 55 -62 60 -57
rect 0 -70 5 -65
rect 9 -130 14 -125
rect 42 -157 47 -152
rect 55 -229 60 -224
rect 0 -237 5 -232
rect 9 -297 14 -292
rect 42 -324 47 -319
rect 56 -394 61 -389
rect 1 -402 6 -397
rect 10 -462 15 -457
rect 43 -489 48 -484
<< metal2 >>
rect 9 131 49 135
rect 0 11 4 94
rect 9 39 13 131
rect 45 119 49 131
rect 45 116 55 119
rect 51 102 55 116
rect 0 7 42 11
rect 9 -33 49 -29
rect 0 -153 4 -70
rect 9 -125 13 -33
rect 45 -45 49 -33
rect 45 -48 55 -45
rect 51 -62 55 -48
rect 0 -157 42 -153
rect 9 -200 49 -196
rect 0 -320 4 -237
rect 9 -292 13 -200
rect 45 -212 49 -200
rect 45 -215 55 -212
rect 51 -229 55 -215
rect 0 -324 42 -320
rect 10 -365 50 -361
rect 1 -485 5 -402
rect 10 -457 14 -365
rect 46 -377 50 -365
rect 46 -380 56 -377
rect 52 -394 56 -380
rect 1 -489 43 -485
<< labels >>
rlabel metal1 26 125 26 125 5 VDD
rlabel metal1 29 80 29 80 1 GND
rlabel metal1 26 65 26 65 5 VDD
rlabel metal1 29 20 29 20 1 GND
rlabel metal1 70 66 70 66 5 VDD
rlabel metal1 84 2 84 2 1 GND
rlabel metal1 70 144 70 144 5 VDD
rlabel metal1 84 80 84 80 1 GND
rlabel metal1 154 109 154 109 5 VDD
rlabel metal1 155 37 155 37 1 GND
rlabel ndcontact 26 89 26 89 1 GND
rlabel pdcontact 26 114 26 114 1 VDD
rlabel ndcontact 57 93 57 93 1 GND
rlabel pdcontact 60 132 60 132 1 VDD
rlabel pdcontact 80 132 80 132 1 VDD
rlabel pdcontact 100 132 100 132 1 VDD
rlabel ndcontact 100 90 100 90 1 GND
rlabel ndcontact 145 46 145 46 1 GND
rlabel ndcontact 165 46 165 46 1 GND
rlabel ndcontact 185 46 185 46 1 GND
rlabel pdcontact 185 71 185 71 1 VDD
rlabel pdcontact 185 -260 185 -260 1 VDD
rlabel ndcontact 185 -285 185 -285 1 GND
rlabel ndcontact 165 -285 165 -285 1 GND
rlabel ndcontact 145 -285 145 -285 1 GND
rlabel ndcontact 100 -319 100 -319 1 GND
rlabel pdcontact 100 -277 100 -277 1 VDD
rlabel ndcontact 100 -241 100 -241 1 GND
rlabel pdcontact 100 -199 100 -199 1 VDD
rlabel pdcontact 80 -199 80 -199 1 VDD
rlabel pdcontact 60 -199 60 -199 1 VDD
rlabel ndcontact 57 -238 57 -238 1 GND
rlabel pdcontact 80 -277 80 -277 1 VDD
rlabel pdcontact 60 -277 60 -277 1 VDD
rlabel ndcontact 57 -316 57 -316 1 GND
rlabel pdcontact 26 -217 26 -217 1 VDD
rlabel ndcontact 26 -242 26 -242 1 GND
rlabel pdcontact 26 -277 26 -277 1 VDD
rlabel ndcontact 26 -302 26 -302 1 GND
rlabel metal1 155 -294 155 -294 1 GND
rlabel metal1 154 -222 154 -222 5 VDD
rlabel metal1 84 -251 84 -251 1 GND
rlabel metal1 70 -187 70 -187 5 VDD
rlabel metal1 84 -329 84 -329 1 GND
rlabel metal1 70 -265 70 -265 5 VDD
rlabel metal1 29 -311 29 -311 1 GND
rlabel metal1 26 -266 26 -266 5 VDD
rlabel metal1 29 -251 29 -251 1 GND
rlabel metal1 26 -206 26 -206 5 VDD
rlabel metal1 26 -39 26 -39 5 VDD
rlabel metal1 29 -84 29 -84 1 GND
rlabel metal1 26 -99 26 -99 5 VDD
rlabel metal1 29 -144 29 -144 1 GND
rlabel metal1 70 -98 70 -98 5 VDD
rlabel metal1 84 -162 84 -162 1 GND
rlabel metal1 70 -20 70 -20 5 VDD
rlabel metal1 84 -84 84 -84 1 GND
rlabel metal1 154 -55 154 -55 5 VDD
rlabel metal1 155 -127 155 -127 1 GND
rlabel ndcontact 26 -135 26 -135 1 GND
rlabel pdcontact 26 -110 26 -110 1 VDD
rlabel ndcontact 26 -75 26 -75 1 GND
rlabel pdcontact 26 -50 26 -50 1 VDD
rlabel ndcontact 57 -149 57 -149 1 GND
rlabel pdcontact 60 -110 60 -110 1 VDD
rlabel pdcontact 80 -110 80 -110 1 VDD
rlabel ndcontact 57 -71 57 -71 1 GND
rlabel pdcontact 60 -32 60 -32 1 VDD
rlabel pdcontact 80 -32 80 -32 1 VDD
rlabel pdcontact 100 -32 100 -32 1 VDD
rlabel ndcontact 100 -74 100 -74 1 GND
rlabel pdcontact 100 -110 100 -110 1 VDD
rlabel ndcontact 100 -152 100 -152 1 GND
rlabel ndcontact 145 -118 145 -118 1 GND
rlabel ndcontact 165 -118 165 -118 1 GND
rlabel ndcontact 185 -118 185 -118 1 GND
rlabel pdcontact 185 -93 185 -93 1 VDD
rlabel metal1 27 -371 27 -371 5 VDD
rlabel metal1 30 -416 30 -416 1 GND
rlabel metal1 27 -431 27 -431 5 VDD
rlabel metal1 30 -476 30 -476 1 GND
rlabel metal1 71 -430 71 -430 5 VDD
rlabel metal1 85 -494 85 -494 1 GND
rlabel metal1 71 -352 71 -352 5 VDD
rlabel metal1 85 -416 85 -416 1 GND
rlabel metal1 155 -387 155 -387 5 VDD
rlabel metal1 156 -459 156 -459 1 GND
rlabel ndcontact 27 -467 27 -467 1 GND
rlabel pdcontact 27 -442 27 -442 1 VDD
rlabel ndcontact 27 -407 27 -407 1 GND
rlabel pdcontact 27 -382 27 -382 1 VDD
rlabel ndcontact 58 -481 58 -481 1 GND
rlabel pdcontact 61 -442 61 -442 1 VDD
rlabel pdcontact 81 -442 81 -442 1 VDD
rlabel ndcontact 58 -403 58 -403 1 GND
rlabel pdcontact 61 -364 61 -364 1 VDD
rlabel pdcontact 81 -364 81 -364 1 VDD
rlabel pdcontact 101 -364 101 -364 1 VDD
rlabel ndcontact 101 -406 101 -406 1 GND
rlabel pdcontact 101 -442 101 -442 1 VDD
rlabel ndcontact 101 -484 101 -484 1 GND
rlabel ndcontact 146 -450 146 -450 1 GND
rlabel ndcontact 166 -450 166 -450 1 GND
rlabel ndcontact 186 -450 186 -450 1 GND
rlabel pdcontact 186 -425 186 -425 1 VDD
rlabel polycontact 27 37 27 37 1 p0
rlabel pdcontact 34 54 34 54 1 p0_bar
rlabel polycontact 61 33 61 33 1 p0_bar
rlabel polycontact 73 26 73 26 1 c0
rlabel polycontact 27 97 27 97 1 c0
rlabel pdcontact 34 114 34 114 1 c0_bar
rlabel polycontact 61 113 61 113 1 c0_bar
rlabel polycontact 73 110 73 110 1 p0
rlabel metal1 197 54 197 54 7 s0
rlabel ndcontact 193 46 193 46 1 s0
rlabel pdcontact 193 71 193 71 1 s0
rlabel pdcontact 145 91 145 91 1 vdd
rlabel pdcontact 70 132 70 132 1 a1n
rlabel ndiffusion 70 93 70 93 1 a1m
rlabel ndcontact 82 93 82 93 1 a1n
rlabel polycontact 104 117 104 117 1 a1n
rlabel ndcontact 114 90 114 90 1 outa1
rlabel pdcontact 114 132 114 132 1 outa1
rlabel polycontact 150 68 150 68 1 outa1
rlabel polycontact 158 61 158 61 1 outa2
rlabel polycontact 186 54 186 54 1 s0_bar
rlabel ndcontact 155 46 155 46 1 s0_bar
rlabel pdcontact 165 91 165 91 1 s0_bar
rlabel pdcontact 114 54 114 54 1 outa2
rlabel ndcontact 114 12 114 12 1 outa2
rlabel polycontact 104 37 104 37 1 a2n
rlabel pdcontact 70 54 70 54 1 a2n
rlabel ndcontact 82 15 82 15 1 a2n
rlabel ndiffusion 70 15 70 15 1 a2m
rlabel polycontact 27 -127 27 -127 1 p1
rlabel ndcontact 34 -135 34 -135 1 p1_bar
rlabel pdcontact 34 -110 34 -110 1 p1_bar
rlabel polycontact 61 -131 61 -131 1 p1_bar
rlabel polycontact 73 -138 73 -138 1 c1
rlabel pdcontact 70 -110 70 -110 1 b2n
rlabel ndcontact 82 -149 82 -149 1 b2n
rlabel ndiffusion 70 -149 70 -149 1 b2m
rlabel polycontact 104 -127 104 -127 1 b2n
rlabel pdcontact 114 -110 114 -110 1 outb2
rlabel ndcontact 114 -152 114 -152 1 outb2
rlabel polycontact 158 -103 158 -103 1 outb2
rlabel ndcontact 155 -118 155 -118 1 s1_bar
rlabel polycontact 186 -110 186 -110 1 s1_bar
rlabel metal1 197 -110 197 -110 7 s1
rlabel ndcontact 193 -118 193 -118 1 s1
rlabel pdcontact 193 -93 193 -93 1 s1
rlabel pdcontact 165 -73 165 -73 1 s1_bar
rlabel pdcontact 145 -73 145 -73 1 vdd
rlabel polycontact 150 -96 150 -96 1 outb1
rlabel ndcontact 114 -74 114 -74 1 outb1
rlabel pdcontact 114 -32 114 -32 1 outb1
rlabel polycontact 104 -47 104 -47 1 b1n
rlabel pdcontact 70 -32 70 -32 1 b1n
rlabel ndcontact 82 -71 82 -71 1 b1n
rlabel ndiffusion 70 -71 70 -71 1 b1m
rlabel polycontact 73 -54 73 -54 1 p1
rlabel polycontact 61 -51 61 -51 1 c1_bar
rlabel ndcontact 34 -75 34 -75 1 c1_bar
rlabel pdcontact 34 -50 34 -50 1 c1_bar
rlabel polycontact 27 -67 27 -67 1 c1
rlabel polycontact 27 -294 27 -294 1 p2
rlabel ndcontact 34 -302 34 -302 1 p2_bar
rlabel pdcontact 34 -277 34 -277 1 p2_bar
rlabel polycontact 61 -298 61 -298 1 p2_bar
rlabel polycontact 73 -305 73 -305 1 c2
rlabel polycontact 27 -234 27 -234 1 c2
rlabel ndcontact 34 -242 34 -242 1 c2_bar
rlabel pdcontact 34 -217 34 -217 1 c2_bar
rlabel polycontact 61 -218 61 -218 1 c2_bar
rlabel polycontact 73 -221 73 -221 1 p2
rlabel pdcontact 70 -199 70 -199 1 c1n
rlabel ndcontact 82 -238 82 -238 1 c1n
rlabel ndiffusion 70 -238 70 -238 1 c1m
rlabel polycontact 104 -214 104 -214 1 c1n
rlabel pdcontact 114 -199 114 -199 1 outc1
rlabel ndcontact 114 -241 114 -241 1 outc1
rlabel polycontact 150 -263 150 -263 1 outc1
rlabel pdcontact 145 -240 145 -240 1 vdd
rlabel polycontact 158 -270 158 -270 1 outc2
rlabel pdcontact 165 -240 165 -240 1 s2_bar
rlabel polycontact 186 -277 186 -277 1 s2_bar
rlabel ndcontact 155 -285 155 -285 1 s2_bar
rlabel metal1 197 -277 197 -277 7 s2
rlabel pdcontact 70 -277 70 -277 1 c2n
rlabel ndiffusion 70 -316 70 -316 1 c2m
rlabel ndcontact 82 -316 82 -316 1 c2n
rlabel polycontact 104 -294 104 -294 1 c2n
rlabel ndcontact 114 -319 114 -319 1 outc2
rlabel pdcontact 114 -277 114 -277 1 outc2
rlabel polycontact 28 -459 28 -459 1 p3
rlabel ndcontact 35 -467 35 -467 1 p3_bar
rlabel pdcontact 35 -442 35 -442 1 p3_bar
rlabel polycontact 62 -463 62 -463 1 p3_bar
rlabel polycontact 74 -470 74 -470 1 c3
rlabel polycontact 28 -399 28 -399 1 c3
rlabel ndcontact 35 -407 35 -407 1 c3_bar
rlabel pdcontact 35 -382 35 -382 1 c3_bar
rlabel polycontact 62 -383 62 -383 1 c3_bar
rlabel polycontact 74 -386 74 -386 1 p3
rlabel pdcontact 71 -364 71 -364 1 d1n
rlabel ndcontact 83 -403 83 -403 1 d1n
rlabel ndiffusion 71 -403 71 -403 1 d1m
rlabel polycontact 105 -379 105 -379 1 d1n
rlabel pdcontact 115 -364 115 -364 1 outd1
rlabel ndcontact 115 -406 115 -406 1 outd1
rlabel polycontact 151 -428 151 -428 1 outd1
rlabel polycontact 159 -435 159 -435 1 outd2
rlabel pdcontact 146 -405 146 -405 1 vdd
rlabel pdcontact 166 -405 166 -405 1 s3_bar
rlabel polycontact 187 -442 187 -442 1 s3_bar
rlabel metal1 198 -442 198 -442 7 s3
rlabel pdcontact 194 -425 194 -425 1 s3
rlabel ndcontact 156 -450 156 -450 1 s3_bar
rlabel pdcontact 71 -442 71 -442 1 d2n
rlabel ndcontact 83 -481 83 -481 1 d2n
rlabel ndiffusion 71 -481 71 -481 1 d2m
rlabel polycontact 105 -459 105 -459 1 d2n
rlabel pdcontact 115 -442 115 -442 1 outd2
rlabel ndcontact 115 -484 115 -484 1 outd2
rlabel pdiffusion 156 -404 156 -404 1 dps
rlabel pdiffusion 155 -240 155 -240 1 cps
rlabel pdiffusion 155 -72 155 -72 1 bps
rlabel pdiffusion 155 90 155 90 1 aps
rlabel ndcontact 193 -285 193 -285 1 s2
rlabel pdcontact 193 -260 193 -260 1 s2
rlabel ndcontact 194 -450 194 -450 1 s3
rlabel ndcontact 34 89 34 89 1 c0_bar
rlabel ndcontact 34 29 34 29 1 p0_bar
rlabel pdcontact 26 54 26 54 1 vdd
rlabel ndcontact 26 29 26 29 1 gnd
rlabel ndcontact 57 15 57 15 1 gnd
rlabel pdcontact 60 54 60 54 1 vdd
rlabel pdcontact 80 54 80 54 1 vdd
rlabel ndcontact 100 12 100 12 1 gnd
rlabel pdcontact 100 54 100 54 1 vdd
<< end >>
