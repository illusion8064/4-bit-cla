magic
tech scmos
timestamp 1732009319
<< nwell >>
rect 18 87 42 111
rect 52 105 122 129
rect 137 70 173 94
rect 137 58 201 70
rect 18 27 42 51
rect 52 27 122 51
rect 177 44 201 58
rect 130 -12 201 12
rect 18 -75 42 -51
rect 52 -57 122 -33
rect 134 -92 170 -68
rect 134 -104 198 -92
rect 18 -135 42 -111
rect 52 -135 122 -111
rect 174 -118 198 -104
rect 127 -174 198 -150
rect 18 -237 42 -213
rect 52 -219 122 -195
rect 137 -254 173 -230
rect 137 -266 201 -254
rect 18 -297 42 -273
rect 52 -297 122 -273
rect 177 -280 201 -266
rect 130 -336 201 -312
rect 18 -399 42 -375
rect 52 -381 122 -357
rect 134 -416 170 -392
rect 134 -428 198 -416
rect 18 -459 42 -435
rect 52 -459 122 -435
rect 174 -442 198 -428
rect 127 -498 198 -474
<< ntransistor >>
rect 29 71 31 77
rect 63 72 65 84
rect 75 72 77 84
rect 106 72 108 78
rect 29 11 31 17
rect 63 -6 65 6
rect 75 -6 77 6
rect 150 28 152 34
rect 158 28 160 34
rect 188 28 190 34
rect 106 -6 108 0
rect 141 -45 143 -33
rect 153 -45 155 -33
rect 184 -45 186 -39
rect 29 -91 31 -85
rect 63 -90 65 -78
rect 75 -90 77 -78
rect 106 -90 108 -84
rect 29 -151 31 -145
rect 63 -168 65 -156
rect 75 -168 77 -156
rect 147 -134 149 -128
rect 155 -134 157 -128
rect 185 -134 187 -128
rect 106 -168 108 -162
rect 138 -207 140 -195
rect 150 -207 152 -195
rect 181 -207 183 -201
rect 29 -253 31 -247
rect 63 -252 65 -240
rect 75 -252 77 -240
rect 106 -252 108 -246
rect 29 -313 31 -307
rect 63 -330 65 -318
rect 75 -330 77 -318
rect 150 -296 152 -290
rect 158 -296 160 -290
rect 188 -296 190 -290
rect 106 -330 108 -324
rect 141 -369 143 -357
rect 153 -369 155 -357
rect 184 -369 186 -363
rect 29 -415 31 -409
rect 63 -414 65 -402
rect 75 -414 77 -402
rect 106 -414 108 -408
rect 29 -475 31 -469
rect 63 -492 65 -480
rect 75 -492 77 -480
rect 147 -458 149 -452
rect 155 -458 157 -452
rect 185 -458 187 -452
rect 106 -492 108 -486
rect 138 -531 140 -519
rect 150 -531 152 -519
rect 181 -531 183 -525
<< ptransistor >>
rect 63 111 65 123
rect 75 111 77 123
rect 106 111 108 123
rect 29 93 31 105
rect 150 64 152 88
rect 158 64 160 88
rect 29 33 31 45
rect 63 33 65 45
rect 75 33 77 45
rect 106 33 108 45
rect 188 50 190 62
rect 141 -6 143 6
rect 153 -6 155 6
rect 184 -6 186 6
rect 63 -51 65 -39
rect 75 -51 77 -39
rect 106 -51 108 -39
rect 29 -69 31 -57
rect 147 -98 149 -74
rect 155 -98 157 -74
rect 29 -129 31 -117
rect 63 -129 65 -117
rect 75 -129 77 -117
rect 106 -129 108 -117
rect 185 -112 187 -100
rect 138 -168 140 -156
rect 150 -168 152 -156
rect 181 -168 183 -156
rect 63 -213 65 -201
rect 75 -213 77 -201
rect 106 -213 108 -201
rect 29 -231 31 -219
rect 150 -260 152 -236
rect 158 -260 160 -236
rect 29 -291 31 -279
rect 63 -291 65 -279
rect 75 -291 77 -279
rect 106 -291 108 -279
rect 188 -274 190 -262
rect 141 -330 143 -318
rect 153 -330 155 -318
rect 184 -330 186 -318
rect 63 -375 65 -363
rect 75 -375 77 -363
rect 106 -375 108 -363
rect 29 -393 31 -381
rect 147 -422 149 -398
rect 155 -422 157 -398
rect 29 -453 31 -441
rect 63 -453 65 -441
rect 75 -453 77 -441
rect 106 -453 108 -441
rect 185 -436 187 -424
rect 138 -492 140 -480
rect 150 -492 152 -480
rect 181 -492 183 -480
<< ndiffusion >>
rect 28 71 29 77
rect 31 71 32 77
rect 59 72 63 84
rect 65 72 75 84
rect 77 72 80 84
rect 102 72 106 78
rect 108 72 112 78
rect 28 11 29 17
rect 31 11 32 17
rect 59 -6 63 6
rect 65 -6 75 6
rect 77 -6 80 6
rect 147 28 150 34
rect 152 28 153 34
rect 157 28 158 34
rect 160 28 163 34
rect 187 28 188 34
rect 190 28 191 34
rect 102 -6 106 0
rect 108 -6 112 0
rect 137 -45 141 -33
rect 143 -45 153 -33
rect 155 -45 158 -33
rect 180 -45 184 -39
rect 186 -45 190 -39
rect 28 -91 29 -85
rect 31 -91 32 -85
rect 59 -90 63 -78
rect 65 -90 75 -78
rect 77 -90 80 -78
rect 102 -90 106 -84
rect 108 -90 112 -84
rect 28 -151 29 -145
rect 31 -151 32 -145
rect 59 -168 63 -156
rect 65 -168 75 -156
rect 77 -168 80 -156
rect 144 -134 147 -128
rect 149 -134 150 -128
rect 154 -134 155 -128
rect 157 -134 160 -128
rect 184 -134 185 -128
rect 187 -134 188 -128
rect 102 -168 106 -162
rect 108 -168 112 -162
rect 134 -207 138 -195
rect 140 -207 150 -195
rect 152 -207 155 -195
rect 177 -207 181 -201
rect 183 -207 187 -201
rect 28 -253 29 -247
rect 31 -253 32 -247
rect 59 -252 63 -240
rect 65 -252 75 -240
rect 77 -252 80 -240
rect 102 -252 106 -246
rect 108 -252 112 -246
rect 28 -313 29 -307
rect 31 -313 32 -307
rect 59 -330 63 -318
rect 65 -330 75 -318
rect 77 -330 80 -318
rect 147 -296 150 -290
rect 152 -296 153 -290
rect 157 -296 158 -290
rect 160 -296 163 -290
rect 187 -296 188 -290
rect 190 -296 191 -290
rect 102 -330 106 -324
rect 108 -330 112 -324
rect 137 -369 141 -357
rect 143 -369 153 -357
rect 155 -369 158 -357
rect 180 -369 184 -363
rect 186 -369 190 -363
rect 28 -415 29 -409
rect 31 -415 32 -409
rect 59 -414 63 -402
rect 65 -414 75 -402
rect 77 -414 80 -402
rect 102 -414 106 -408
rect 108 -414 112 -408
rect 28 -475 29 -469
rect 31 -475 32 -469
rect 59 -492 63 -480
rect 65 -492 75 -480
rect 77 -492 80 -480
rect 144 -458 147 -452
rect 149 -458 150 -452
rect 154 -458 155 -452
rect 157 -458 160 -452
rect 184 -458 185 -452
rect 187 -458 188 -452
rect 102 -492 106 -486
rect 108 -492 112 -486
rect 134 -531 138 -519
rect 140 -531 150 -519
rect 152 -531 155 -519
rect 177 -531 181 -525
rect 183 -531 187 -525
<< pdiffusion >>
rect 62 111 63 123
rect 65 111 68 123
rect 72 111 75 123
rect 77 111 78 123
rect 102 111 106 123
rect 108 111 112 123
rect 28 93 29 105
rect 31 93 32 105
rect 147 64 150 88
rect 152 64 158 88
rect 160 64 163 88
rect 28 33 29 45
rect 31 33 32 45
rect 62 33 63 45
rect 65 33 68 45
rect 72 33 75 45
rect 77 33 78 45
rect 102 33 106 45
rect 108 33 112 45
rect 187 50 188 62
rect 190 50 191 62
rect 140 -6 141 6
rect 143 -6 146 6
rect 150 -6 153 6
rect 155 -6 156 6
rect 180 -6 184 6
rect 186 -6 190 6
rect 62 -51 63 -39
rect 65 -51 68 -39
rect 72 -51 75 -39
rect 77 -51 78 -39
rect 102 -51 106 -39
rect 108 -51 112 -39
rect 28 -69 29 -57
rect 31 -69 32 -57
rect 144 -98 147 -74
rect 149 -98 155 -74
rect 157 -98 160 -74
rect 28 -129 29 -117
rect 31 -129 32 -117
rect 62 -129 63 -117
rect 65 -129 68 -117
rect 72 -129 75 -117
rect 77 -129 78 -117
rect 102 -129 106 -117
rect 108 -129 112 -117
rect 184 -112 185 -100
rect 187 -112 188 -100
rect 137 -168 138 -156
rect 140 -168 143 -156
rect 147 -168 150 -156
rect 152 -168 153 -156
rect 177 -168 181 -156
rect 183 -168 187 -156
rect 62 -213 63 -201
rect 65 -213 68 -201
rect 72 -213 75 -201
rect 77 -213 78 -201
rect 102 -213 106 -201
rect 108 -213 112 -201
rect 28 -231 29 -219
rect 31 -231 32 -219
rect 147 -260 150 -236
rect 152 -260 158 -236
rect 160 -260 163 -236
rect 28 -291 29 -279
rect 31 -291 32 -279
rect 62 -291 63 -279
rect 65 -291 68 -279
rect 72 -291 75 -279
rect 77 -291 78 -279
rect 102 -291 106 -279
rect 108 -291 112 -279
rect 187 -274 188 -262
rect 190 -274 191 -262
rect 140 -330 141 -318
rect 143 -330 146 -318
rect 150 -330 153 -318
rect 155 -330 156 -318
rect 180 -330 184 -318
rect 186 -330 190 -318
rect 62 -375 63 -363
rect 65 -375 68 -363
rect 72 -375 75 -363
rect 77 -375 78 -363
rect 102 -375 106 -363
rect 108 -375 112 -363
rect 28 -393 29 -381
rect 31 -393 32 -381
rect 144 -422 147 -398
rect 149 -422 155 -398
rect 157 -422 160 -398
rect 28 -453 29 -441
rect 31 -453 32 -441
rect 62 -453 63 -441
rect 65 -453 68 -441
rect 72 -453 75 -441
rect 77 -453 78 -441
rect 102 -453 106 -441
rect 108 -453 112 -441
rect 184 -436 185 -424
rect 187 -436 188 -424
rect 137 -492 138 -480
rect 140 -492 143 -480
rect 147 -492 150 -480
rect 152 -492 153 -480
rect 177 -492 181 -480
rect 183 -492 187 -480
<< ndcontact >>
rect 24 71 28 77
rect 32 71 36 77
rect 55 72 59 84
rect 80 72 84 84
rect 98 72 102 78
rect 112 72 116 78
rect 24 11 28 17
rect 32 11 36 17
rect 55 -6 59 6
rect 80 -6 84 6
rect 143 28 147 34
rect 153 28 157 34
rect 163 28 167 34
rect 183 28 187 34
rect 191 28 195 34
rect 98 -6 102 0
rect 112 -6 116 0
rect 133 -45 137 -33
rect 158 -45 162 -33
rect 176 -45 180 -39
rect 190 -45 194 -39
rect 24 -91 28 -85
rect 32 -91 36 -85
rect 55 -90 59 -78
rect 80 -90 84 -78
rect 98 -90 102 -84
rect 112 -90 116 -84
rect 24 -151 28 -145
rect 32 -151 36 -145
rect 55 -168 59 -156
rect 80 -168 84 -156
rect 140 -134 144 -128
rect 150 -134 154 -128
rect 160 -134 164 -128
rect 180 -134 184 -128
rect 188 -134 192 -128
rect 98 -168 102 -162
rect 112 -168 116 -162
rect 130 -207 134 -195
rect 155 -207 159 -195
rect 173 -207 177 -201
rect 187 -207 191 -201
rect 24 -253 28 -247
rect 32 -253 36 -247
rect 55 -252 59 -240
rect 80 -252 84 -240
rect 98 -252 102 -246
rect 112 -252 116 -246
rect 24 -313 28 -307
rect 32 -313 36 -307
rect 55 -330 59 -318
rect 80 -330 84 -318
rect 143 -296 147 -290
rect 153 -296 157 -290
rect 163 -296 167 -290
rect 183 -296 187 -290
rect 191 -296 195 -290
rect 98 -330 102 -324
rect 112 -330 116 -324
rect 133 -369 137 -357
rect 158 -369 162 -357
rect 176 -369 180 -363
rect 190 -369 194 -363
rect 24 -415 28 -409
rect 32 -415 36 -409
rect 55 -414 59 -402
rect 80 -414 84 -402
rect 98 -414 102 -408
rect 112 -414 116 -408
rect 24 -475 28 -469
rect 32 -475 36 -469
rect 55 -492 59 -480
rect 80 -492 84 -480
rect 140 -458 144 -452
rect 150 -458 154 -452
rect 160 -458 164 -452
rect 180 -458 184 -452
rect 188 -458 192 -452
rect 98 -492 102 -486
rect 112 -492 116 -486
rect 130 -531 134 -519
rect 155 -531 159 -519
rect 173 -531 177 -525
rect 187 -531 191 -525
<< pdcontact >>
rect 58 111 62 123
rect 68 111 72 123
rect 78 111 82 123
rect 98 111 102 123
rect 112 111 116 123
rect 24 93 28 105
rect 32 93 36 105
rect 143 64 147 88
rect 163 64 167 88
rect 24 33 28 45
rect 32 33 36 45
rect 58 33 62 45
rect 68 33 72 45
rect 78 33 82 45
rect 98 33 102 45
rect 112 33 116 45
rect 183 50 187 62
rect 191 50 195 62
rect 136 -6 140 6
rect 146 -6 150 6
rect 156 -6 160 6
rect 176 -6 180 6
rect 190 -6 194 6
rect 58 -51 62 -39
rect 68 -51 72 -39
rect 78 -51 82 -39
rect 98 -51 102 -39
rect 112 -51 116 -39
rect 24 -69 28 -57
rect 32 -69 36 -57
rect 140 -98 144 -74
rect 160 -98 164 -74
rect 24 -129 28 -117
rect 32 -129 36 -117
rect 58 -129 62 -117
rect 68 -129 72 -117
rect 78 -129 82 -117
rect 98 -129 102 -117
rect 112 -129 116 -117
rect 180 -112 184 -100
rect 188 -112 192 -100
rect 133 -168 137 -156
rect 143 -168 147 -156
rect 153 -168 157 -156
rect 173 -168 177 -156
rect 187 -168 191 -156
rect 58 -213 62 -201
rect 68 -213 72 -201
rect 78 -213 82 -201
rect 98 -213 102 -201
rect 112 -213 116 -201
rect 24 -231 28 -219
rect 32 -231 36 -219
rect 143 -260 147 -236
rect 163 -260 167 -236
rect 24 -291 28 -279
rect 32 -291 36 -279
rect 58 -291 62 -279
rect 68 -291 72 -279
rect 78 -291 82 -279
rect 98 -291 102 -279
rect 112 -291 116 -279
rect 183 -274 187 -262
rect 191 -274 195 -262
rect 136 -330 140 -318
rect 146 -330 150 -318
rect 156 -330 160 -318
rect 176 -330 180 -318
rect 190 -330 194 -318
rect 58 -375 62 -363
rect 68 -375 72 -363
rect 78 -375 82 -363
rect 98 -375 102 -363
rect 112 -375 116 -363
rect 24 -393 28 -381
rect 32 -393 36 -381
rect 140 -422 144 -398
rect 160 -422 164 -398
rect 24 -453 28 -441
rect 32 -453 36 -441
rect 58 -453 62 -441
rect 68 -453 72 -441
rect 78 -453 82 -441
rect 98 -453 102 -441
rect 112 -453 116 -441
rect 180 -436 184 -424
rect 188 -436 192 -424
rect 133 -492 137 -480
rect 143 -492 147 -480
rect 153 -492 157 -480
rect 173 -492 177 -480
rect 187 -492 191 -480
<< polysilicon >>
rect 63 123 65 126
rect 75 123 77 126
rect 106 123 108 126
rect 29 105 31 108
rect 29 77 31 93
rect 63 84 65 111
rect 75 84 77 111
rect 106 78 108 111
rect 150 88 152 91
rect 158 88 160 91
rect 29 68 31 71
rect 63 69 65 72
rect 75 69 77 72
rect 106 69 108 72
rect 150 55 152 64
rect 29 45 31 48
rect 63 45 65 48
rect 75 45 77 48
rect 106 45 108 48
rect 150 34 152 51
rect 158 48 160 64
rect 188 62 190 65
rect 158 34 160 44
rect 188 34 190 50
rect 29 17 31 33
rect 29 8 31 11
rect 63 6 65 33
rect 75 6 77 33
rect 106 0 108 33
rect 150 25 152 28
rect 158 25 160 28
rect 188 24 190 28
rect 141 6 143 9
rect 153 6 155 9
rect 184 6 186 9
rect 63 -9 65 -6
rect 75 -9 77 -6
rect 106 -9 108 -6
rect 141 -33 143 -6
rect 153 -33 155 -6
rect 63 -39 65 -36
rect 75 -39 77 -36
rect 106 -39 108 -36
rect 184 -39 186 -6
rect 141 -48 143 -45
rect 153 -48 155 -45
rect 184 -48 186 -45
rect 29 -57 31 -54
rect 29 -85 31 -69
rect 63 -78 65 -51
rect 75 -78 77 -51
rect 106 -84 108 -51
rect 147 -74 149 -71
rect 155 -74 157 -71
rect 29 -94 31 -91
rect 63 -93 65 -90
rect 75 -93 77 -90
rect 106 -93 108 -90
rect 147 -107 149 -98
rect 29 -117 31 -114
rect 63 -117 65 -114
rect 75 -117 77 -114
rect 106 -117 108 -114
rect 147 -128 149 -111
rect 155 -114 157 -98
rect 185 -100 187 -97
rect 155 -128 157 -118
rect 185 -128 187 -112
rect 29 -145 31 -129
rect 29 -154 31 -151
rect 63 -156 65 -129
rect 75 -156 77 -129
rect 106 -162 108 -129
rect 147 -137 149 -134
rect 155 -137 157 -134
rect 185 -138 187 -134
rect 138 -156 140 -153
rect 150 -156 152 -153
rect 181 -156 183 -153
rect 63 -171 65 -168
rect 75 -171 77 -168
rect 106 -171 108 -168
rect 138 -195 140 -168
rect 150 -195 152 -168
rect 63 -201 65 -198
rect 75 -201 77 -198
rect 106 -201 108 -198
rect 181 -201 183 -168
rect 138 -210 140 -207
rect 150 -210 152 -207
rect 181 -210 183 -207
rect 29 -219 31 -216
rect 29 -247 31 -231
rect 63 -240 65 -213
rect 75 -240 77 -213
rect 106 -246 108 -213
rect 150 -236 152 -233
rect 158 -236 160 -233
rect 29 -256 31 -253
rect 63 -255 65 -252
rect 75 -255 77 -252
rect 106 -255 108 -252
rect 150 -269 152 -260
rect 29 -279 31 -276
rect 63 -279 65 -276
rect 75 -279 77 -276
rect 106 -279 108 -276
rect 150 -290 152 -273
rect 158 -276 160 -260
rect 188 -262 190 -259
rect 158 -290 160 -280
rect 188 -290 190 -274
rect 29 -307 31 -291
rect 29 -316 31 -313
rect 63 -318 65 -291
rect 75 -318 77 -291
rect 106 -324 108 -291
rect 150 -299 152 -296
rect 158 -299 160 -296
rect 188 -300 190 -296
rect 141 -318 143 -315
rect 153 -318 155 -315
rect 184 -318 186 -315
rect 63 -333 65 -330
rect 75 -333 77 -330
rect 106 -333 108 -330
rect 141 -357 143 -330
rect 153 -357 155 -330
rect 63 -363 65 -360
rect 75 -363 77 -360
rect 106 -363 108 -360
rect 184 -363 186 -330
rect 141 -372 143 -369
rect 153 -372 155 -369
rect 184 -372 186 -369
rect 29 -381 31 -378
rect 29 -409 31 -393
rect 63 -402 65 -375
rect 75 -402 77 -375
rect 106 -408 108 -375
rect 147 -398 149 -395
rect 155 -398 157 -395
rect 29 -418 31 -415
rect 63 -417 65 -414
rect 75 -417 77 -414
rect 106 -417 108 -414
rect 147 -431 149 -422
rect 29 -441 31 -438
rect 63 -441 65 -438
rect 75 -441 77 -438
rect 106 -441 108 -438
rect 147 -452 149 -435
rect 155 -438 157 -422
rect 185 -424 187 -421
rect 155 -452 157 -442
rect 185 -452 187 -436
rect 29 -469 31 -453
rect 29 -478 31 -475
rect 63 -480 65 -453
rect 75 -480 77 -453
rect 106 -486 108 -453
rect 147 -461 149 -458
rect 155 -461 157 -458
rect 185 -462 187 -458
rect 138 -480 140 -477
rect 150 -480 152 -477
rect 181 -480 183 -477
rect 63 -495 65 -492
rect 75 -495 77 -492
rect 106 -495 108 -492
rect 138 -519 140 -492
rect 150 -519 152 -492
rect 181 -525 183 -492
rect 138 -534 140 -531
rect 150 -534 152 -531
rect 181 -534 183 -531
<< polycontact >>
rect 59 96 63 100
rect 25 80 29 84
rect 71 93 75 97
rect 102 100 106 104
rect 148 51 152 55
rect 156 44 160 48
rect 184 37 188 41
rect 25 20 29 24
rect 59 16 63 20
rect 71 9 75 13
rect 102 20 106 24
rect 137 -23 141 -19
rect 149 -30 153 -26
rect 180 -19 184 -15
rect 59 -66 63 -62
rect 25 -82 29 -78
rect 71 -69 75 -65
rect 102 -62 106 -58
rect 145 -111 149 -107
rect 153 -118 157 -114
rect 181 -125 185 -121
rect 25 -142 29 -138
rect 59 -146 63 -142
rect 71 -153 75 -149
rect 102 -142 106 -138
rect 134 -185 138 -181
rect 146 -192 150 -188
rect 177 -181 181 -177
rect 59 -228 63 -224
rect 25 -244 29 -240
rect 71 -231 75 -227
rect 102 -224 106 -220
rect 148 -273 152 -269
rect 156 -280 160 -276
rect 184 -287 188 -283
rect 25 -304 29 -300
rect 59 -308 63 -304
rect 71 -315 75 -311
rect 102 -304 106 -300
rect 137 -347 141 -343
rect 149 -354 153 -350
rect 180 -343 184 -339
rect 59 -390 63 -386
rect 25 -406 29 -402
rect 71 -393 75 -389
rect 102 -386 106 -382
rect 145 -435 149 -431
rect 153 -442 157 -438
rect 181 -449 185 -445
rect 25 -466 29 -462
rect 59 -470 63 -466
rect 71 -477 75 -473
rect 102 -466 106 -462
rect 134 -509 138 -505
rect 146 -516 150 -512
rect 177 -505 181 -501
<< metal1 >>
rect 52 127 102 131
rect 58 123 62 127
rect 78 123 82 127
rect 18 109 42 113
rect 98 123 102 127
rect 24 105 28 109
rect 68 104 72 111
rect 68 100 102 104
rect 112 102 116 111
rect 32 84 36 93
rect 46 96 59 100
rect 46 84 50 96
rect 67 91 71 97
rect 60 87 71 91
rect 80 84 84 100
rect 5 80 25 84
rect 32 80 50 84
rect 32 77 36 80
rect 112 98 134 102
rect 112 78 116 98
rect 24 67 28 71
rect 55 67 59 72
rect 98 67 102 72
rect 18 63 42 67
rect 52 63 102 67
rect 130 55 134 98
rect 137 92 176 96
rect 143 88 147 92
rect 172 70 176 92
rect 172 66 187 70
rect 18 49 42 53
rect 52 49 102 53
rect 130 51 148 55
rect 24 45 28 49
rect 58 45 62 49
rect 78 45 82 49
rect 98 45 102 49
rect 32 24 36 33
rect 68 24 72 33
rect 112 24 116 33
rect 130 44 156 48
rect 130 24 134 44
rect 163 41 167 64
rect 183 62 187 66
rect 191 41 195 50
rect 153 37 184 41
rect 191 37 199 41
rect 153 34 157 37
rect 191 34 195 37
rect 143 24 147 28
rect 163 24 167 28
rect 183 24 187 28
rect 14 20 25 24
rect 32 20 54 24
rect 68 20 102 24
rect 112 20 134 24
rect 137 20 187 24
rect 32 17 36 20
rect 50 16 59 20
rect 24 7 28 11
rect 47 9 71 13
rect 18 3 42 7
rect 9 -17 13 2
rect 47 -8 51 9
rect 80 6 84 20
rect 112 0 116 20
rect 130 10 180 14
rect 136 6 140 10
rect 156 6 160 10
rect 176 6 180 10
rect 55 -11 59 -6
rect 98 -11 102 -6
rect 52 -14 102 -11
rect 146 -15 150 -6
rect 190 -15 194 -6
rect 9 -19 117 -17
rect 146 -19 180 -15
rect 190 -19 198 -15
rect 9 -21 137 -19
rect 113 -23 137 -21
rect 5 -26 110 -24
rect 5 -28 149 -26
rect 106 -30 149 -28
rect 52 -35 102 -31
rect 158 -33 162 -19
rect 58 -39 62 -35
rect 78 -39 82 -35
rect 18 -53 42 -49
rect 98 -39 102 -35
rect 190 -39 194 -19
rect 133 -50 137 -45
rect 176 -50 180 -45
rect 24 -57 28 -53
rect 68 -58 72 -51
rect 68 -62 102 -58
rect 112 -60 116 -51
rect 130 -54 180 -50
rect 32 -78 36 -69
rect 46 -66 59 -62
rect 46 -78 50 -66
rect 67 -71 71 -65
rect 60 -75 71 -71
rect 80 -78 84 -62
rect 5 -82 25 -78
rect 32 -82 50 -78
rect 32 -85 36 -82
rect 112 -64 131 -60
rect 112 -84 116 -64
rect 24 -95 28 -91
rect 55 -95 59 -90
rect 98 -95 102 -90
rect 18 -99 42 -95
rect 52 -99 102 -95
rect 127 -107 131 -64
rect 134 -70 173 -66
rect 140 -74 144 -70
rect 169 -92 173 -70
rect 169 -96 184 -92
rect 18 -113 42 -109
rect 52 -113 102 -109
rect 127 -111 145 -107
rect 24 -117 28 -113
rect 58 -117 62 -113
rect 78 -117 82 -113
rect 98 -117 102 -113
rect 32 -138 36 -129
rect 68 -138 72 -129
rect 112 -138 116 -129
rect 127 -118 153 -114
rect 127 -138 131 -118
rect 160 -121 164 -98
rect 180 -100 184 -96
rect 188 -121 192 -112
rect 150 -125 181 -121
rect 188 -125 196 -121
rect 150 -128 154 -125
rect 188 -128 192 -125
rect 140 -138 144 -134
rect 160 -138 164 -134
rect 180 -138 184 -134
rect 14 -142 25 -138
rect 32 -142 54 -138
rect 68 -142 102 -138
rect 112 -142 131 -138
rect 134 -142 184 -138
rect 32 -145 36 -142
rect 50 -146 59 -142
rect 24 -155 28 -151
rect 47 -153 71 -149
rect 18 -159 42 -155
rect 9 -179 13 -160
rect 47 -170 51 -153
rect 80 -156 84 -142
rect 112 -162 116 -142
rect 127 -152 177 -148
rect 133 -156 137 -152
rect 153 -156 157 -152
rect 173 -156 177 -152
rect 55 -173 59 -168
rect 98 -173 102 -168
rect 52 -176 102 -173
rect 143 -177 147 -168
rect 187 -177 191 -168
rect 9 -181 117 -179
rect 143 -181 177 -177
rect 187 -181 195 -177
rect 9 -183 134 -181
rect 113 -185 134 -183
rect 5 -188 110 -186
rect 5 -190 146 -188
rect 106 -192 146 -190
rect 52 -197 102 -193
rect 155 -195 159 -181
rect 58 -201 62 -197
rect 78 -201 82 -197
rect 18 -215 42 -211
rect 98 -201 102 -197
rect 187 -201 191 -181
rect 130 -212 134 -207
rect 173 -212 177 -207
rect 24 -219 28 -215
rect 68 -220 72 -213
rect 68 -224 102 -220
rect 112 -222 116 -213
rect 127 -216 177 -212
rect 32 -240 36 -231
rect 46 -228 59 -224
rect 46 -240 50 -228
rect 67 -233 71 -227
rect 60 -237 71 -233
rect 80 -240 84 -224
rect 5 -244 25 -240
rect 32 -244 50 -240
rect 32 -247 36 -244
rect 112 -226 134 -222
rect 112 -246 116 -226
rect 24 -257 28 -253
rect 55 -257 59 -252
rect 98 -257 102 -252
rect 18 -261 42 -257
rect 52 -261 102 -257
rect 130 -269 134 -226
rect 137 -232 176 -228
rect 143 -236 147 -232
rect 172 -254 176 -232
rect 172 -258 187 -254
rect 18 -275 42 -271
rect 52 -275 102 -271
rect 130 -273 148 -269
rect 24 -279 28 -275
rect 58 -279 62 -275
rect 78 -279 82 -275
rect 98 -279 102 -275
rect 32 -300 36 -291
rect 68 -300 72 -291
rect 112 -300 116 -291
rect 130 -280 156 -276
rect 130 -300 134 -280
rect 163 -283 167 -260
rect 183 -262 187 -258
rect 191 -283 195 -274
rect 153 -287 184 -283
rect 191 -287 199 -283
rect 153 -290 157 -287
rect 191 -290 195 -287
rect 143 -300 147 -296
rect 163 -300 167 -296
rect 183 -300 187 -296
rect 14 -304 25 -300
rect 32 -304 54 -300
rect 68 -304 102 -300
rect 112 -304 134 -300
rect 137 -304 187 -300
rect 32 -307 36 -304
rect 50 -308 59 -304
rect 24 -317 28 -313
rect 47 -315 71 -311
rect 18 -321 42 -317
rect 9 -341 13 -322
rect 47 -332 51 -315
rect 80 -318 84 -304
rect 112 -324 116 -304
rect 130 -314 180 -310
rect 136 -318 140 -314
rect 156 -318 160 -314
rect 176 -318 180 -314
rect 55 -335 59 -330
rect 98 -335 102 -330
rect 52 -338 102 -335
rect 146 -339 150 -330
rect 190 -339 194 -330
rect 9 -343 117 -341
rect 146 -343 180 -339
rect 190 -343 198 -339
rect 9 -345 137 -343
rect 113 -347 137 -345
rect 5 -350 110 -348
rect 5 -352 149 -350
rect 106 -354 149 -352
rect 52 -359 102 -355
rect 158 -357 162 -343
rect 58 -363 62 -359
rect 78 -363 82 -359
rect 18 -377 42 -373
rect 98 -363 102 -359
rect 190 -363 194 -343
rect 133 -374 137 -369
rect 176 -374 180 -369
rect 24 -381 28 -377
rect 68 -382 72 -375
rect 68 -386 102 -382
rect 112 -384 116 -375
rect 130 -378 180 -374
rect 32 -402 36 -393
rect 46 -390 59 -386
rect 46 -402 50 -390
rect 67 -395 71 -389
rect 60 -399 71 -395
rect 80 -402 84 -386
rect 5 -406 25 -402
rect 32 -406 50 -402
rect 32 -409 36 -406
rect 112 -388 131 -384
rect 112 -408 116 -388
rect 24 -419 28 -415
rect 55 -419 59 -414
rect 98 -419 102 -414
rect 18 -423 42 -419
rect 52 -423 102 -419
rect 127 -431 131 -388
rect 134 -394 173 -390
rect 140 -398 144 -394
rect 169 -416 173 -394
rect 169 -420 184 -416
rect 18 -437 42 -433
rect 52 -437 102 -433
rect 127 -435 145 -431
rect 24 -441 28 -437
rect 58 -441 62 -437
rect 78 -441 82 -437
rect 98 -441 102 -437
rect 32 -462 36 -453
rect 68 -462 72 -453
rect 112 -462 116 -453
rect 127 -442 153 -438
rect 127 -462 131 -442
rect 160 -445 164 -422
rect 180 -424 184 -420
rect 188 -445 192 -436
rect 150 -449 181 -445
rect 188 -449 196 -445
rect 150 -452 154 -449
rect 188 -452 192 -449
rect 140 -462 144 -458
rect 160 -462 164 -458
rect 180 -462 184 -458
rect 14 -466 25 -462
rect 32 -466 54 -462
rect 68 -466 102 -462
rect 112 -466 131 -462
rect 134 -466 184 -462
rect 32 -469 36 -466
rect 50 -470 59 -466
rect 24 -479 28 -475
rect 47 -477 71 -473
rect 18 -483 42 -479
rect 9 -503 13 -484
rect 47 -494 51 -477
rect 80 -480 84 -466
rect 112 -486 116 -466
rect 127 -476 177 -472
rect 133 -480 137 -476
rect 153 -480 157 -476
rect 173 -480 177 -476
rect 55 -497 59 -492
rect 98 -497 102 -492
rect 52 -500 102 -497
rect 143 -501 147 -492
rect 187 -501 191 -492
rect 9 -505 117 -503
rect 143 -505 177 -501
rect 187 -505 195 -501
rect 9 -507 134 -505
rect 113 -509 134 -507
rect 5 -512 110 -510
rect 5 -514 146 -512
rect 106 -516 146 -514
rect 155 -519 159 -505
rect 187 -525 191 -505
rect 130 -536 134 -531
rect 173 -536 177 -531
rect 127 -540 177 -536
<< m2contact >>
rect 55 87 60 92
rect 0 79 5 84
rect 9 19 14 24
rect 9 2 14 7
rect 42 -8 47 -3
rect 0 -28 5 -23
rect 55 -75 60 -70
rect 0 -83 5 -78
rect 9 -143 14 -138
rect 9 -160 14 -155
rect 42 -170 47 -165
rect 0 -190 5 -185
rect 55 -237 60 -232
rect 0 -245 5 -240
rect 9 -305 14 -300
rect 9 -322 14 -317
rect 42 -332 47 -327
rect 0 -352 5 -347
rect 55 -399 60 -394
rect 0 -407 5 -402
rect 9 -467 14 -462
rect 9 -484 14 -479
rect 42 -494 47 -489
rect 0 -514 5 -509
<< metal2 >>
rect 9 116 49 120
rect 0 -4 4 79
rect 9 24 13 116
rect 45 104 49 116
rect 45 101 55 104
rect 51 87 55 101
rect 9 7 13 19
rect 0 -8 42 -4
rect 0 -23 4 -8
rect 9 -46 49 -42
rect 0 -166 4 -83
rect 9 -138 13 -46
rect 45 -58 49 -46
rect 45 -61 55 -58
rect 51 -75 55 -61
rect 9 -155 13 -143
rect 0 -170 42 -166
rect 0 -185 4 -170
rect 9 -208 49 -204
rect 0 -328 4 -245
rect 9 -300 13 -208
rect 45 -220 49 -208
rect 45 -223 55 -220
rect 51 -237 55 -223
rect 9 -317 13 -305
rect 0 -332 42 -328
rect 0 -347 4 -332
rect 9 -370 49 -366
rect 0 -490 4 -407
rect 9 -462 13 -370
rect 45 -382 49 -370
rect 45 -385 55 -382
rect 51 -399 55 -385
rect 9 -479 13 -467
rect 0 -494 42 -490
rect 0 -509 4 -494
<< labels >>
rlabel metal1 26 110 26 110 5 VDD
rlabel metal1 29 65 29 65 1 GND
rlabel metal1 26 50 26 50 5 VDD
rlabel metal1 29 5 29 5 1 GND
rlabel metal1 70 51 70 51 5 VDD
rlabel metal1 84 -13 84 -13 1 GND
rlabel metal1 70 129 70 129 5 VDD
rlabel metal1 84 65 84 65 1 GND
rlabel metal1 154 94 154 94 5 VDD
rlabel metal1 155 22 155 22 1 GND
rlabel ndcontact 26 14 26 14 1 GND
rlabel pdcontact 26 39 26 39 1 VDD
rlabel ndcontact 26 74 26 74 1 GND
rlabel pdcontact 26 99 26 99 1 VDD
rlabel ndcontact 57 0 57 0 1 GND
rlabel ndiffusion 70 0 70 0 1 and2m
rlabel ndcontact 82 0 82 0 1 and2n
rlabel pdcontact 60 39 60 39 1 VDD
rlabel pdcontact 70 39 70 39 1 and2n
rlabel pdcontact 80 39 80 39 1 VDD
rlabel ndcontact 57 78 57 78 1 GND
rlabel ndiffusion 70 78 70 78 1 and1m
rlabel ndcontact 82 78 82 78 1 and1n
rlabel pdcontact 60 117 60 117 1 VDD
rlabel pdcontact 80 117 80 117 1 VDD
rlabel pdcontact 70 117 70 117 1 and1n
rlabel polycontact 104 102 104 102 1 and1n
rlabel pdcontact 100 117 100 117 1 VDD
rlabel pdcontact 114 117 114 117 1 outand1
rlabel ndcontact 114 75 114 75 1 outand1
rlabel ndcontact 100 75 100 75 1 GND
rlabel pdcontact 100 39 100 39 1 VDD
rlabel pdcontact 114 39 114 39 1 outand2
rlabel ndcontact 114 -3 114 -3 1 outand2
rlabel ndcontact 100 -3 100 -3 1 GND
rlabel polycontact 104 22 104 22 1 and2n
rlabel polycontact 150 53 150 53 1 outand1
rlabel polycontact 158 46 158 46 1 outand2
rlabel ndcontact 145 31 145 31 1 GND
rlabel ndcontact 165 31 165 31 1 GND
rlabel ndcontact 185 31 185 31 1 GND
rlabel pdcontact 185 56 185 56 1 VDD
rlabel metal1 135 -52 135 -52 2 GND
rlabel metal1 148 12 148 12 5 VDD
rlabel metal1 26 -52 26 -52 5 VDD
rlabel metal1 29 -97 29 -97 1 GND
rlabel metal1 26 -112 26 -112 5 VDD
rlabel metal1 29 -157 29 -157 1 GND
rlabel metal1 70 -111 70 -111 5 VDD
rlabel metal1 84 -175 84 -175 1 GND
rlabel metal1 70 -33 70 -33 5 VDD
rlabel metal1 84 -97 84 -97 1 GND
rlabel ndcontact 26 -148 26 -148 1 GND
rlabel pdcontact 26 -123 26 -123 1 VDD
rlabel ndcontact 26 -88 26 -88 1 GND
rlabel pdcontact 26 -63 26 -63 1 VDD
rlabel ndcontact 57 -162 57 -162 1 GND
rlabel pdcontact 60 -123 60 -123 1 VDD
rlabel pdcontact 80 -123 80 -123 1 VDD
rlabel ndcontact 57 -84 57 -84 1 GND
rlabel pdcontact 60 -45 60 -45 1 VDD
rlabel pdcontact 80 -45 80 -45 1 VDD
rlabel pdcontact 100 -45 100 -45 1 VDD
rlabel ndcontact 100 -87 100 -87 1 GND
rlabel pdcontact 100 -123 100 -123 1 VDD
rlabel ndcontact 100 -165 100 -165 1 GND
rlabel metal1 151 -68 151 -68 5 VDD
rlabel metal1 152 -140 152 -140 1 GND
rlabel ndcontact 142 -131 142 -131 1 GND
rlabel ndcontact 162 -131 162 -131 1 GND
rlabel ndcontact 182 -131 182 -131 1 GND
rlabel pdcontact 182 -106 182 -106 1 VDD
rlabel metal1 145 -150 145 -150 5 VDD
rlabel metal1 132 -214 132 -214 2 GND
rlabel metal1 26 -214 26 -214 5 VDD
rlabel metal1 29 -259 29 -259 1 GND
rlabel metal1 26 -274 26 -274 5 VDD
rlabel metal1 29 -319 29 -319 1 GND
rlabel metal1 70 -273 70 -273 5 VDD
rlabel metal1 84 -337 84 -337 1 GND
rlabel metal1 70 -195 70 -195 5 VDD
rlabel metal1 84 -259 84 -259 1 GND
rlabel metal1 154 -230 154 -230 5 VDD
rlabel metal1 155 -302 155 -302 1 GND
rlabel ndcontact 26 -310 26 -310 1 GND
rlabel pdcontact 26 -285 26 -285 1 VDD
rlabel ndcontact 26 -250 26 -250 1 GND
rlabel pdcontact 26 -225 26 -225 1 VDD
rlabel ndcontact 57 -324 57 -324 1 GND
rlabel pdcontact 60 -285 60 -285 1 VDD
rlabel pdcontact 80 -285 80 -285 1 VDD
rlabel ndcontact 57 -246 57 -246 1 GND
rlabel pdcontact 60 -207 60 -207 1 VDD
rlabel pdcontact 80 -207 80 -207 1 VDD
rlabel pdcontact 100 -207 100 -207 1 VDD
rlabel ndcontact 100 -249 100 -249 1 GND
rlabel pdcontact 100 -285 100 -285 1 VDD
rlabel ndcontact 100 -327 100 -327 1 GND
rlabel ndcontact 145 -293 145 -293 1 GND
rlabel ndcontact 165 -293 165 -293 1 GND
rlabel ndcontact 185 -293 185 -293 1 GND
rlabel pdcontact 185 -268 185 -268 1 VDD
rlabel metal1 135 -376 135 -376 2 GND
rlabel metal1 148 -312 148 -312 5 VDD
rlabel metal1 26 -376 26 -376 5 VDD
rlabel metal1 29 -421 29 -421 1 GND
rlabel metal1 26 -436 26 -436 5 VDD
rlabel metal1 29 -481 29 -481 1 GND
rlabel metal1 70 -435 70 -435 5 VDD
rlabel metal1 84 -499 84 -499 1 GND
rlabel metal1 70 -357 70 -357 5 VDD
rlabel metal1 84 -421 84 -421 1 GND
rlabel ndcontact 26 -472 26 -472 1 GND
rlabel pdcontact 26 -447 26 -447 1 VDD
rlabel ndcontact 26 -412 26 -412 1 GND
rlabel pdcontact 26 -387 26 -387 1 VDD
rlabel ndcontact 57 -486 57 -486 1 GND
rlabel pdcontact 60 -447 60 -447 1 VDD
rlabel pdcontact 80 -447 80 -447 1 VDD
rlabel ndcontact 57 -408 57 -408 1 GND
rlabel pdcontact 60 -369 60 -369 1 VDD
rlabel pdcontact 80 -369 80 -369 1 VDD
rlabel pdcontact 100 -369 100 -369 1 VDD
rlabel ndcontact 100 -411 100 -411 1 GND
rlabel pdcontact 100 -447 100 -447 1 VDD
rlabel ndcontact 100 -489 100 -489 1 GND
rlabel metal1 151 -392 151 -392 5 VDD
rlabel metal1 152 -464 152 -464 1 GND
rlabel ndcontact 142 -455 142 -455 1 GND
rlabel ndcontact 162 -455 162 -455 1 GND
rlabel ndcontact 182 -455 182 -455 1 GND
rlabel pdcontact 182 -430 182 -430 1 VDD
rlabel metal1 145 -474 145 -474 5 VDD
rlabel metal1 132 -538 132 -538 2 GND
rlabel metal1 196 -17 196 -17 7 g0
rlabel ndcontact 192 -42 192 -42 1 g0
rlabel pdcontact 192 0 192 0 1 g0
rlabel ndcontact 178 -42 178 -42 1 gnd
rlabel ndcontact 160 -39 160 -39 1 g0_bar
rlabel polycontact 182 -17 182 -17 1 g0_bar
rlabel pdcontact 148 0 148 0 1 g0_bar
rlabel pdcontact 178 0 178 0 1 vdd
rlabel pdcontact 158 0 158 0 1 vdd
rlabel pdcontact 138 0 138 0 1 vdd
rlabel ndcontact 135 -39 135 -39 1 gnd
rlabel ndiffusion 147 -39 147 -39 1 and0m
rlabel polycontact 151 -28 151 -28 1 b0
rlabel ndcontact 193 31 193 31 1 p0
rlabel metal1 197 39 197 39 7 p0
rlabel pdcontact 193 56 193 56 1 p0
rlabel polycontact 186 39 186 39 1 p0_bar
rlabel ndcontact 155 31 155 31 1 p0_bar
rlabel pdcontact 165 76 165 76 1 p0_bar
rlabel pdcontact 145 76 145 76 1 vdd
rlabel polycontact 27 22 27 22 1 a0
rlabel ndcontact 34 14 34 14 1 a0_bar
rlabel pdcontact 34 39 34 39 1 a0_bar
rlabel polycontact 61 18 61 18 1 a0_bar
rlabel polycontact 73 11 73 11 1 b0
rlabel polycontact 27 82 27 82 1 b0
rlabel pdcontact 34 99 34 99 1 b0_bar
rlabel ndcontact 34 74 34 74 1 b0_bar
rlabel polycontact 61 98 61 98 1 b0_bar
rlabel polycontact 73 95 73 95 1 a0
rlabel polycontact 139 -21 139 -21 1 a0
rlabel ndcontact 175 -204 175 -204 1 gnd
rlabel ndcontact 189 -204 189 -204 1 g1
rlabel metal1 193 -179 193 -179 1 g1
rlabel pdcontact 189 -162 189 -162 1 g1
rlabel pdcontact 175 -162 175 -162 1 vdd
rlabel polycontact 179 -179 179 -179 1 g1_bar
rlabel ndcontact 157 -201 157 -201 1 g1_bar
rlabel ndcontact 132 -201 132 -201 1 gnd
rlabel pdcontact 145 -162 145 -162 1 g1_bar
rlabel pdcontact 155 -162 155 -162 1 vdd
rlabel pdcontact 135 -162 135 -162 1 vdd
rlabel polycontact 148 -190 148 -190 1 b1
rlabel polycontact 136 -183 136 -183 1 a1
rlabel metal1 194 -123 194 -123 1 p1
rlabel ndcontact 190 -131 190 -131 1 p1
rlabel pdcontact 190 -106 190 -106 1 p1
rlabel polycontact 183 -123 183 -123 1 p1_bar
rlabel ndcontact 152 -131 152 -131 1 p1_bar
rlabel pdcontact 162 -86 162 -86 1 p1_bar
rlabel pdcontact 142 -86 142 -86 1 vdd
rlabel polycontact 27 -140 27 -140 1 a1
rlabel ndcontact 34 -148 34 -148 1 a1_bar
rlabel pdcontact 34 -123 34 -123 1 a1_bar
rlabel polycontact 61 -144 61 -144 1 a1_bar
rlabel polycontact 73 -151 73 -151 1 b1
rlabel polycontact 27 -80 27 -80 1 b1
rlabel ndcontact 34 -88 34 -88 1 b1_bar
rlabel pdcontact 34 -63 34 -63 1 b1_bar
rlabel polycontact 61 -64 61 -64 1 b1_bar
rlabel polycontact 73 -67 73 -67 1 a1
rlabel metal1 196 -341 196 -341 7 g2
rlabel ndcontact 192 -366 192 -366 1 g2
rlabel pdcontact 192 -324 192 -324 1 g2
rlabel ndcontact 178 -366 178 -366 1 gnd
rlabel ndcontact 160 -363 160 -363 1 g2_bar
rlabel ndcontact 135 -363 135 -363 1 gnd
rlabel polycontact 182 -341 182 -341 1 g2_bar
rlabel polycontact 151 -352 151 -352 1 b2
rlabel polycontact 139 -345 139 -345 1 a2
rlabel pdcontact 178 -324 178 -324 1 vdd
rlabel pdcontact 158 -324 158 -324 1 vdd
rlabel pdcontact 138 -324 138 -324 1 vdd
rlabel pdcontact 148 -324 148 -324 1 g2_bar
rlabel ndcontact 193 -293 193 -293 1 p2
rlabel metal1 197 -285 197 -285 7 p2
rlabel pdcontact 193 -268 193 -268 1 p2
rlabel polycontact 186 -285 186 -285 1 p2_bar
rlabel ndcontact 155 -293 155 -293 1 p2_bar
rlabel pdcontact 165 -249 165 -249 1 p2_bar
rlabel pdcontact 145 -248 145 -248 1 vdd
rlabel polycontact 27 -302 27 -302 1 a2
rlabel ndcontact 34 -310 34 -310 1 a2_bar
rlabel pdcontact 34 -285 34 -285 1 a2_bar
rlabel polycontact 61 -306 61 -306 1 a2_bar
rlabel polycontact 73 -313 73 -313 1 b2
rlabel polycontact 27 -242 27 -242 1 b2
rlabel pdcontact 34 -225 34 -225 1 b2_bar
rlabel ndcontact 34 -250 34 -250 1 b2_bar
rlabel polycontact 61 -226 61 -226 1 b2_bar
rlabel polycontact 73 -229 73 -229 1 a2
rlabel ndcontact 175 -528 175 -528 1 gnd
rlabel ndcontact 189 -528 189 -528 1 g3
rlabel metal1 193 -503 193 -503 1 g3
rlabel pdcontact 189 -486 189 -486 1 g3
rlabel pdcontact 175 -486 175 -486 1 vdd
rlabel polycontact 179 -503 179 -503 1 g3_bar
rlabel ndcontact 157 -525 157 -525 1 g3_bar
rlabel ndcontact 132 -525 132 -525 1 gnd
rlabel polycontact 148 -514 148 -514 1 b3
rlabel polycontact 136 -507 136 -507 1 a3
rlabel pdcontact 155 -486 155 -486 1 vdd
rlabel pdcontact 135 -486 135 -486 1 vdd
rlabel pdcontact 145 -486 145 -486 1 g3_bar
rlabel ndcontact 190 -455 190 -455 1 p3
rlabel metal1 194 -447 194 -447 1 p3
rlabel pdcontact 190 -430 190 -430 1 p3
rlabel polycontact 183 -447 183 -447 1 p3_bar
rlabel ndcontact 152 -455 152 -455 1 p3_bar
rlabel pdcontact 162 -410 162 -410 1 p3_bar
rlabel pdcontact 142 -410 142 -410 1 vdd
rlabel polycontact 27 -464 27 -464 1 a3
rlabel ndcontact 34 -472 34 -472 1 a3_bar
rlabel pdcontact 34 -447 34 -447 1 a3_bar
rlabel polycontact 61 -468 61 -468 1 a3_bar
rlabel polycontact 73 -475 73 -475 1 b3
rlabel polycontact 27 -404 27 -404 1 b3
rlabel pdcontact 34 -387 34 -387 1 b3_bar
rlabel ndcontact 34 -412 34 -412 1 b3_bar
rlabel polycontact 61 -388 61 -388 1 b3_bar
rlabel polycontact 73 -391 73 -391 1 a3
rlabel pdcontact 70 -45 70 -45 1 anda1n
rlabel ndcontact 82 -84 82 -84 1 anda1n
rlabel ndiffusion 70 -84 70 -84 1 anda1m
rlabel polycontact 104 -60 104 -60 1 anda1n
rlabel pdcontact 114 -45 114 -45 1 outanda1
rlabel ndcontact 114 -87 114 -87 1 outanda1
rlabel polycontact 147 -109 147 -109 1 outanda1
rlabel polycontact 155 -116 155 -116 1 outanda2
rlabel pdcontact 114 -123 114 -123 1 outanda2
rlabel ndcontact 114 -165 114 -165 1 outanda2
rlabel polycontact 104 -140 104 -140 1 anda2n
rlabel ndcontact 82 -162 82 -162 1 anda2n
rlabel ndiffusion 70 -162 70 -162 1 anda2m
rlabel pdcontact 70 -123 70 -123 1 anda2n
rlabel pdcontact 70 -207 70 -207 1 andb1n
rlabel ndiffusion 70 -246 70 -246 1 andb1m
rlabel ndcontact 82 -246 82 -246 1 andb1n
rlabel polycontact 104 -222 104 -222 1 andb1n
rlabel pdcontact 114 -207 114 -207 1 outband1
rlabel ndcontact 114 -249 114 -249 1 outband1
rlabel polycontact 150 -271 150 -271 1 outband1
rlabel polycontact 158 -278 158 -278 1 outband2
rlabel pdcontact 114 -285 114 -285 1 outband2
rlabel ndcontact 114 -327 114 -327 1 outband2
rlabel polycontact 104 -302 104 -302 1 andb2n
rlabel pdcontact 70 -285 70 -285 1 andb2n
rlabel ndcontact 82 -324 82 -324 1 andb2n
rlabel ndiffusion 70 -324 70 -324 1 andb2m
rlabel pdcontact 70 -369 70 -369 1 andc1n
rlabel ndcontact 82 -408 82 -408 1 andc1n
rlabel ndiffusion 70 -408 70 -408 1 andc1m
rlabel polycontact 104 -384 104 -384 1 andc1n
rlabel pdcontact 114 -369 114 -369 1 outcand1
rlabel ndcontact 114 -411 114 -411 1 outcand1
rlabel polycontact 147 -433 147 -433 1 outcand1
rlabel polycontact 155 -440 155 -440 1 outcand2
rlabel pdcontact 114 -447 114 -447 1 outcand2
rlabel ndcontact 114 -489 114 -489 1 outcand2
rlabel polycontact 104 -464 104 -464 1 andc2n
rlabel ndcontact 82 -486 82 -486 1 andc2n
rlabel ndiffusion 70 -486 70 -486 1 andc2m
rlabel pdcontact 70 -447 70 -447 1 andc2n
<< end >>
