magic
tech scmos
timestamp 1732041806
<< nwell >>
rect -215 -234 -80 -210
rect -215 -246 -175 -234
rect -215 -341 -80 -317
rect -215 -353 -175 -341
rect 10 -385 34 -361
rect 44 -367 114 -343
rect 129 -402 165 -378
rect 529 -400 553 -376
rect 563 -382 633 -358
rect 129 -414 193 -402
rect -215 -448 -80 -424
rect 10 -445 34 -421
rect 44 -445 114 -421
rect 169 -428 193 -414
rect 648 -417 684 -393
rect -215 -460 -175 -448
rect 290 -452 360 -428
rect 370 -452 406 -428
rect 648 -429 712 -417
rect 122 -484 193 -460
rect 370 -464 434 -452
rect 529 -460 553 -436
rect 563 -460 633 -436
rect 688 -443 712 -429
rect 410 -478 434 -464
rect 780 -465 915 -441
rect 780 -477 820 -465
rect -215 -555 -80 -531
rect 10 -547 34 -523
rect 44 -529 114 -505
rect 290 -539 371 -515
rect -215 -567 -175 -555
rect 126 -564 162 -540
rect 387 -556 431 -546
rect 126 -576 190 -564
rect 10 -607 34 -583
rect 44 -607 114 -583
rect 166 -590 190 -576
rect 387 -582 460 -556
rect 529 -564 553 -540
rect 563 -546 633 -522
rect 648 -581 684 -557
rect 780 -572 915 -548
rect 648 -593 712 -581
rect 780 -584 820 -572
rect -215 -662 -80 -638
rect 119 -646 190 -622
rect 290 -634 360 -610
rect 529 -624 553 -600
rect 563 -624 633 -600
rect 688 -607 712 -593
rect -215 -674 -175 -662
rect 10 -709 34 -685
rect 44 -691 114 -667
rect 780 -679 915 -655
rect 129 -726 165 -702
rect 290 -723 378 -699
rect 129 -738 193 -726
rect -215 -769 -80 -745
rect 10 -769 34 -745
rect 44 -769 114 -745
rect 169 -752 193 -738
rect 387 -747 439 -730
rect 529 -731 553 -707
rect 563 -713 633 -689
rect 780 -691 820 -679
rect 387 -766 474 -747
rect 648 -748 684 -724
rect 648 -760 712 -748
rect -215 -781 -175 -769
rect 442 -773 474 -766
rect 122 -808 193 -784
rect 529 -791 553 -767
rect 563 -791 633 -767
rect 688 -774 712 -760
rect 780 -786 915 -762
rect 290 -821 371 -797
rect 780 -798 820 -786
rect -215 -876 -80 -852
rect 10 -871 34 -847
rect 44 -853 114 -829
rect -215 -888 -175 -876
rect 126 -888 162 -864
rect 126 -900 190 -888
rect 10 -931 34 -907
rect 44 -931 114 -907
rect 166 -914 190 -900
rect 290 -914 360 -890
rect 530 -896 554 -872
rect 564 -878 634 -854
rect 649 -913 685 -889
rect 780 -893 915 -869
rect 780 -905 820 -893
rect 649 -925 713 -913
rect -215 -983 -80 -959
rect 119 -970 190 -946
rect 530 -956 554 -932
rect 564 -956 634 -932
rect 689 -939 713 -925
rect -215 -995 -175 -983
rect -215 -1090 -80 -1066
rect -215 -1102 -175 -1090
<< ntransistor >>
rect -202 -284 -200 -278
rect -164 -284 -162 -272
rect -152 -284 -150 -272
rect -127 -284 -125 -272
rect -115 -284 -113 -272
rect -93 -284 -91 -278
rect -202 -391 -200 -385
rect -164 -391 -162 -379
rect -152 -391 -150 -379
rect -127 -391 -125 -379
rect -115 -391 -113 -379
rect -93 -391 -91 -385
rect 21 -401 23 -395
rect 55 -400 57 -388
rect 67 -400 69 -388
rect 98 -400 100 -394
rect 540 -416 542 -410
rect 574 -415 576 -403
rect 586 -415 588 -403
rect 617 -415 619 -409
rect -202 -498 -200 -492
rect -164 -498 -162 -486
rect -152 -498 -150 -486
rect -127 -498 -125 -486
rect -115 -498 -113 -486
rect 21 -461 23 -455
rect 55 -478 57 -466
rect 67 -478 69 -466
rect 142 -444 144 -438
rect 150 -444 152 -438
rect 180 -444 182 -438
rect 98 -478 100 -472
rect -93 -498 -91 -492
rect 133 -517 135 -505
rect 145 -517 147 -505
rect 301 -485 303 -473
rect 313 -485 315 -473
rect 344 -485 346 -479
rect 540 -476 542 -470
rect 383 -494 385 -488
rect 391 -494 393 -488
rect 421 -494 423 -488
rect 574 -493 576 -481
rect 586 -493 588 -481
rect 661 -459 663 -453
rect 669 -459 671 -453
rect 699 -459 701 -453
rect 617 -493 619 -487
rect 176 -517 178 -511
rect 793 -515 795 -509
rect 831 -515 833 -503
rect 843 -515 845 -503
rect 868 -515 870 -503
rect 880 -515 882 -503
rect 902 -515 904 -509
rect -202 -605 -200 -599
rect -164 -605 -162 -593
rect -152 -605 -150 -593
rect -127 -605 -125 -593
rect -115 -605 -113 -593
rect 21 -563 23 -557
rect 55 -562 57 -550
rect 67 -562 69 -550
rect 98 -562 100 -556
rect -93 -605 -91 -599
rect 301 -579 303 -567
rect 313 -579 315 -567
rect 325 -579 327 -567
rect 355 -576 357 -570
rect 21 -623 23 -617
rect 55 -640 57 -628
rect 67 -640 69 -628
rect 139 -606 141 -600
rect 147 -606 149 -600
rect 177 -606 179 -600
rect 540 -580 542 -574
rect 574 -579 576 -567
rect 586 -579 588 -567
rect 617 -579 619 -573
rect 447 -598 449 -592
rect 400 -619 402 -613
rect 408 -619 410 -613
rect 416 -619 418 -613
rect 98 -640 100 -634
rect -202 -712 -200 -706
rect -164 -712 -162 -700
rect -152 -712 -150 -700
rect -127 -712 -125 -700
rect -115 -712 -113 -700
rect 130 -679 132 -667
rect 142 -679 144 -667
rect 301 -667 303 -655
rect 313 -667 315 -655
rect 540 -640 542 -634
rect 574 -657 576 -645
rect 586 -657 588 -645
rect 661 -623 663 -617
rect 669 -623 671 -617
rect 699 -623 701 -617
rect 793 -622 795 -616
rect 831 -622 833 -610
rect 843 -622 845 -610
rect 868 -622 870 -610
rect 880 -622 882 -610
rect 902 -622 904 -616
rect 617 -657 619 -651
rect 344 -667 346 -661
rect 173 -679 175 -673
rect -93 -712 -91 -706
rect 21 -725 23 -719
rect 55 -724 57 -712
rect 67 -724 69 -712
rect 98 -724 100 -718
rect -202 -819 -200 -813
rect -164 -819 -162 -807
rect -152 -819 -150 -807
rect -127 -819 -125 -807
rect -115 -819 -113 -807
rect 21 -785 23 -779
rect 55 -802 57 -790
rect 67 -802 69 -790
rect 142 -768 144 -762
rect 150 -768 152 -762
rect 180 -768 182 -762
rect 301 -770 303 -758
rect 313 -770 315 -758
rect 325 -770 327 -758
rect 337 -770 339 -758
rect 540 -747 542 -741
rect 574 -746 576 -734
rect 586 -746 588 -734
rect 793 -729 795 -723
rect 831 -729 833 -717
rect 843 -729 845 -717
rect 868 -729 870 -717
rect 880 -729 882 -717
rect 902 -729 904 -723
rect 617 -746 619 -740
rect 362 -767 364 -761
rect 98 -802 100 -796
rect -93 -819 -91 -813
rect 133 -841 135 -829
rect 145 -841 147 -829
rect 461 -789 463 -783
rect 400 -811 402 -805
rect 408 -811 410 -805
rect 416 -811 418 -805
rect 424 -811 426 -805
rect 540 -807 542 -801
rect 176 -841 178 -835
rect -202 -926 -200 -920
rect -164 -926 -162 -914
rect -152 -926 -150 -914
rect -127 -926 -125 -914
rect -115 -926 -113 -914
rect 21 -887 23 -881
rect 55 -886 57 -874
rect 67 -886 69 -874
rect 301 -861 303 -849
rect 313 -861 315 -849
rect 325 -861 327 -849
rect 574 -824 576 -812
rect 586 -824 588 -812
rect 661 -790 663 -784
rect 669 -790 671 -784
rect 699 -790 701 -784
rect 617 -824 619 -818
rect 793 -836 795 -830
rect 831 -836 833 -824
rect 843 -836 845 -824
rect 868 -836 870 -824
rect 880 -836 882 -824
rect 902 -836 904 -830
rect 355 -858 357 -852
rect 98 -886 100 -880
rect -93 -926 -91 -920
rect 21 -947 23 -941
rect 55 -964 57 -952
rect 67 -964 69 -952
rect 139 -930 141 -924
rect 147 -930 149 -924
rect 177 -930 179 -924
rect 301 -947 303 -935
rect 313 -947 315 -935
rect 541 -912 543 -906
rect 575 -911 577 -899
rect 587 -911 589 -899
rect 618 -911 620 -905
rect 344 -947 346 -941
rect 793 -943 795 -937
rect 831 -943 833 -931
rect 843 -943 845 -931
rect 868 -943 870 -931
rect 880 -943 882 -931
rect 902 -943 904 -937
rect 98 -964 100 -958
rect -202 -1033 -200 -1027
rect -164 -1033 -162 -1021
rect -152 -1033 -150 -1021
rect -127 -1033 -125 -1021
rect -115 -1033 -113 -1021
rect 130 -1003 132 -991
rect 142 -1003 144 -991
rect 541 -972 543 -966
rect 575 -989 577 -977
rect 587 -989 589 -977
rect 662 -955 664 -949
rect 670 -955 672 -949
rect 700 -955 702 -949
rect 618 -989 620 -983
rect 173 -1003 175 -997
rect -93 -1033 -91 -1027
rect -202 -1140 -200 -1134
rect -164 -1140 -162 -1128
rect -152 -1140 -150 -1128
rect -127 -1140 -125 -1128
rect -115 -1140 -113 -1128
rect -93 -1140 -91 -1134
<< ptransistor >>
rect -202 -240 -200 -216
rect -190 -240 -188 -216
rect -164 -228 -162 -216
rect -127 -228 -125 -216
rect -93 -228 -91 -216
rect -202 -347 -200 -323
rect -190 -347 -188 -323
rect -164 -335 -162 -323
rect -127 -335 -125 -323
rect -93 -335 -91 -323
rect 55 -361 57 -349
rect 67 -361 69 -349
rect 98 -361 100 -349
rect 21 -379 23 -367
rect 574 -376 576 -364
rect 586 -376 588 -364
rect 617 -376 619 -364
rect 142 -408 144 -384
rect 150 -408 152 -384
rect 540 -394 542 -382
rect -202 -454 -200 -430
rect -190 -454 -188 -430
rect -164 -442 -162 -430
rect -127 -442 -125 -430
rect -93 -442 -91 -430
rect 21 -439 23 -427
rect 55 -439 57 -427
rect 67 -439 69 -427
rect 98 -439 100 -427
rect 180 -422 182 -410
rect 661 -423 663 -399
rect 669 -423 671 -399
rect 301 -446 303 -434
rect 313 -446 315 -434
rect 344 -446 346 -434
rect 133 -478 135 -466
rect 145 -478 147 -466
rect 176 -478 178 -466
rect 55 -523 57 -511
rect 67 -523 69 -511
rect 98 -523 100 -511
rect 383 -458 385 -434
rect 391 -458 393 -434
rect 540 -454 542 -442
rect 574 -454 576 -442
rect 586 -454 588 -442
rect 617 -454 619 -442
rect 699 -437 701 -425
rect 421 -472 423 -460
rect 793 -471 795 -447
rect 805 -471 807 -447
rect 831 -459 833 -447
rect 868 -459 870 -447
rect 902 -459 904 -447
rect -202 -561 -200 -537
rect -190 -561 -188 -537
rect -164 -549 -162 -537
rect -127 -549 -125 -537
rect -93 -549 -91 -537
rect 21 -541 23 -529
rect 301 -533 303 -521
rect 313 -533 315 -521
rect 325 -533 327 -521
rect 355 -533 357 -521
rect 139 -570 141 -546
rect 147 -570 149 -546
rect 21 -601 23 -589
rect 55 -601 57 -589
rect 67 -601 69 -589
rect 98 -601 100 -589
rect 177 -584 179 -572
rect 574 -540 576 -528
rect 586 -540 588 -528
rect 617 -540 619 -528
rect 400 -576 402 -552
rect 408 -576 410 -552
rect 416 -576 418 -552
rect 540 -558 542 -546
rect 447 -576 449 -564
rect 661 -587 663 -563
rect 669 -587 671 -563
rect 793 -578 795 -554
rect 805 -578 807 -554
rect 831 -566 833 -554
rect 868 -566 870 -554
rect 902 -566 904 -554
rect 301 -628 303 -616
rect 313 -628 315 -616
rect 344 -628 346 -616
rect 540 -618 542 -606
rect 574 -618 576 -606
rect 586 -618 588 -606
rect 617 -618 619 -606
rect 699 -601 701 -589
rect 130 -640 132 -628
rect 142 -640 144 -628
rect 173 -640 175 -628
rect -202 -668 -200 -644
rect -190 -668 -188 -644
rect -164 -656 -162 -644
rect -127 -656 -125 -644
rect -93 -656 -91 -644
rect 55 -685 57 -673
rect 67 -685 69 -673
rect 98 -685 100 -673
rect 793 -685 795 -661
rect 805 -685 807 -661
rect 831 -673 833 -661
rect 868 -673 870 -661
rect 902 -673 904 -661
rect 21 -703 23 -691
rect 142 -732 144 -708
rect 150 -732 152 -708
rect 301 -717 303 -705
rect 313 -717 315 -705
rect 325 -717 327 -705
rect 337 -717 339 -705
rect 362 -717 364 -705
rect 574 -707 576 -695
rect 586 -707 588 -695
rect 617 -707 619 -695
rect -202 -775 -200 -751
rect -190 -775 -188 -751
rect -164 -763 -162 -751
rect -127 -763 -125 -751
rect -93 -763 -91 -751
rect 21 -763 23 -751
rect 55 -763 57 -751
rect 67 -763 69 -751
rect 98 -763 100 -751
rect 180 -746 182 -734
rect 540 -725 542 -713
rect 400 -760 402 -736
rect 408 -760 410 -736
rect 416 -760 418 -736
rect 424 -760 426 -736
rect 661 -754 663 -730
rect 669 -754 671 -730
rect 133 -802 135 -790
rect 145 -802 147 -790
rect 176 -802 178 -790
rect 55 -847 57 -835
rect 67 -847 69 -835
rect 98 -847 100 -835
rect 301 -815 303 -803
rect 313 -815 315 -803
rect 325 -815 327 -803
rect 355 -815 357 -803
rect 461 -767 463 -755
rect 540 -785 542 -773
rect 574 -785 576 -773
rect 586 -785 588 -773
rect 617 -785 619 -773
rect 699 -768 701 -756
rect -202 -882 -200 -858
rect -190 -882 -188 -858
rect -164 -870 -162 -858
rect -127 -870 -125 -858
rect -93 -870 -91 -858
rect 21 -865 23 -853
rect 793 -792 795 -768
rect 805 -792 807 -768
rect 831 -780 833 -768
rect 868 -780 870 -768
rect 902 -780 904 -768
rect 139 -894 141 -870
rect 147 -894 149 -870
rect 575 -872 577 -860
rect 587 -872 589 -860
rect 618 -872 620 -860
rect 541 -890 543 -878
rect 21 -925 23 -913
rect 55 -925 57 -913
rect 67 -925 69 -913
rect 98 -925 100 -913
rect 177 -908 179 -896
rect 301 -908 303 -896
rect 313 -908 315 -896
rect 344 -908 346 -896
rect 662 -919 664 -895
rect 670 -919 672 -895
rect 793 -899 795 -875
rect 805 -899 807 -875
rect 831 -887 833 -875
rect 868 -887 870 -875
rect 902 -887 904 -875
rect 541 -950 543 -938
rect 575 -950 577 -938
rect 587 -950 589 -938
rect 618 -950 620 -938
rect 700 -933 702 -921
rect 130 -964 132 -952
rect 142 -964 144 -952
rect 173 -964 175 -952
rect -202 -989 -200 -965
rect -190 -989 -188 -965
rect -164 -977 -162 -965
rect -127 -977 -125 -965
rect -93 -977 -91 -965
rect -202 -1096 -200 -1072
rect -190 -1096 -188 -1072
rect -164 -1084 -162 -1072
rect -127 -1084 -125 -1072
rect -93 -1084 -91 -1072
<< ndiffusion >>
rect -205 -284 -202 -278
rect -200 -284 -185 -278
rect -167 -284 -164 -272
rect -162 -284 -152 -272
rect -150 -284 -147 -272
rect -130 -284 -127 -272
rect -125 -284 -115 -272
rect -113 -284 -110 -272
rect -94 -284 -93 -278
rect -91 -284 -90 -278
rect -205 -391 -202 -385
rect -200 -391 -185 -385
rect -167 -391 -164 -379
rect -162 -391 -152 -379
rect -150 -391 -147 -379
rect -130 -391 -127 -379
rect -125 -391 -115 -379
rect -113 -391 -110 -379
rect -94 -391 -93 -385
rect -91 -391 -90 -385
rect 20 -401 21 -395
rect 23 -401 24 -395
rect 51 -400 55 -388
rect 57 -400 67 -388
rect 69 -400 72 -388
rect 94 -400 98 -394
rect 100 -400 104 -394
rect 539 -416 540 -410
rect 542 -416 543 -410
rect 570 -415 574 -403
rect 576 -415 586 -403
rect 588 -415 591 -403
rect 613 -415 617 -409
rect 619 -415 623 -409
rect -205 -498 -202 -492
rect -200 -498 -185 -492
rect -167 -498 -164 -486
rect -162 -498 -152 -486
rect -150 -498 -147 -486
rect -130 -498 -127 -486
rect -125 -498 -115 -486
rect -113 -498 -110 -486
rect 20 -461 21 -455
rect 23 -461 24 -455
rect 51 -478 55 -466
rect 57 -478 67 -466
rect 69 -478 72 -466
rect 139 -444 142 -438
rect 144 -444 145 -438
rect 149 -444 150 -438
rect 152 -444 155 -438
rect 179 -444 180 -438
rect 182 -444 183 -438
rect 94 -478 98 -472
rect 100 -478 104 -472
rect -94 -498 -93 -492
rect -91 -498 -90 -492
rect 129 -517 133 -505
rect 135 -517 145 -505
rect 147 -517 150 -505
rect 297 -485 301 -473
rect 303 -485 313 -473
rect 315 -485 318 -473
rect 340 -485 344 -479
rect 346 -485 350 -479
rect 539 -476 540 -470
rect 542 -476 543 -470
rect 380 -494 383 -488
rect 385 -494 386 -488
rect 390 -494 391 -488
rect 393 -494 396 -488
rect 420 -494 421 -488
rect 423 -494 424 -488
rect 570 -493 574 -481
rect 576 -493 586 -481
rect 588 -493 591 -481
rect 658 -459 661 -453
rect 663 -459 664 -453
rect 668 -459 669 -453
rect 671 -459 674 -453
rect 698 -459 699 -453
rect 701 -459 702 -453
rect 613 -493 617 -487
rect 619 -493 623 -487
rect 172 -517 176 -511
rect 178 -517 182 -511
rect 790 -515 793 -509
rect 795 -515 810 -509
rect 828 -515 831 -503
rect 833 -515 843 -503
rect 845 -515 848 -503
rect 865 -515 868 -503
rect 870 -515 880 -503
rect 882 -515 885 -503
rect 901 -515 902 -509
rect 904 -515 905 -509
rect -205 -605 -202 -599
rect -200 -605 -185 -599
rect -167 -605 -164 -593
rect -162 -605 -152 -593
rect -150 -605 -147 -593
rect -130 -605 -127 -593
rect -125 -605 -115 -593
rect -113 -605 -110 -593
rect 20 -563 21 -557
rect 23 -563 24 -557
rect 51 -562 55 -550
rect 57 -562 67 -550
rect 69 -562 72 -550
rect 94 -562 98 -556
rect 100 -562 104 -556
rect -94 -605 -93 -599
rect -91 -605 -90 -599
rect 297 -579 301 -567
rect 303 -579 313 -567
rect 315 -579 325 -567
rect 327 -579 328 -567
rect 351 -576 355 -570
rect 357 -576 361 -570
rect 20 -623 21 -617
rect 23 -623 24 -617
rect 51 -640 55 -628
rect 57 -640 67 -628
rect 69 -640 72 -628
rect 136 -606 139 -600
rect 141 -606 142 -600
rect 146 -606 147 -600
rect 149 -606 152 -600
rect 176 -606 177 -600
rect 179 -606 180 -600
rect 539 -580 540 -574
rect 542 -580 543 -574
rect 570 -579 574 -567
rect 576 -579 586 -567
rect 588 -579 591 -567
rect 613 -579 617 -573
rect 619 -579 623 -573
rect 446 -598 447 -592
rect 449 -598 450 -592
rect 397 -619 400 -613
rect 402 -619 403 -613
rect 407 -619 408 -613
rect 410 -619 411 -613
rect 415 -619 416 -613
rect 418 -619 421 -613
rect 94 -640 98 -634
rect 100 -640 104 -634
rect -205 -712 -202 -706
rect -200 -712 -185 -706
rect -167 -712 -164 -700
rect -162 -712 -152 -700
rect -150 -712 -147 -700
rect -130 -712 -127 -700
rect -125 -712 -115 -700
rect -113 -712 -110 -700
rect 126 -679 130 -667
rect 132 -679 142 -667
rect 144 -679 147 -667
rect 297 -667 301 -655
rect 303 -667 313 -655
rect 315 -667 318 -655
rect 539 -640 540 -634
rect 542 -640 543 -634
rect 570 -657 574 -645
rect 576 -657 586 -645
rect 588 -657 591 -645
rect 658 -623 661 -617
rect 663 -623 664 -617
rect 668 -623 669 -617
rect 671 -623 674 -617
rect 698 -623 699 -617
rect 701 -623 702 -617
rect 790 -622 793 -616
rect 795 -622 810 -616
rect 828 -622 831 -610
rect 833 -622 843 -610
rect 845 -622 848 -610
rect 865 -622 868 -610
rect 870 -622 880 -610
rect 882 -622 885 -610
rect 901 -622 902 -616
rect 904 -622 905 -616
rect 613 -657 617 -651
rect 619 -657 623 -651
rect 340 -667 344 -661
rect 346 -667 350 -661
rect 169 -679 173 -673
rect 175 -679 179 -673
rect -94 -712 -93 -706
rect -91 -712 -90 -706
rect 20 -725 21 -719
rect 23 -725 24 -719
rect 51 -724 55 -712
rect 57 -724 67 -712
rect 69 -724 72 -712
rect 94 -724 98 -718
rect 100 -724 104 -718
rect -205 -819 -202 -813
rect -200 -819 -185 -813
rect -167 -819 -164 -807
rect -162 -819 -152 -807
rect -150 -819 -147 -807
rect -130 -819 -127 -807
rect -125 -819 -115 -807
rect -113 -819 -110 -807
rect 20 -785 21 -779
rect 23 -785 24 -779
rect 51 -802 55 -790
rect 57 -802 67 -790
rect 69 -802 72 -790
rect 139 -768 142 -762
rect 144 -768 145 -762
rect 149 -768 150 -762
rect 152 -768 155 -762
rect 179 -768 180 -762
rect 182 -768 183 -762
rect 297 -770 301 -758
rect 303 -770 313 -758
rect 315 -770 325 -758
rect 327 -770 337 -758
rect 339 -770 340 -758
rect 539 -747 540 -741
rect 542 -747 543 -741
rect 570 -746 574 -734
rect 576 -746 586 -734
rect 588 -746 591 -734
rect 790 -729 793 -723
rect 795 -729 810 -723
rect 828 -729 831 -717
rect 833 -729 843 -717
rect 845 -729 848 -717
rect 865 -729 868 -717
rect 870 -729 880 -717
rect 882 -729 885 -717
rect 901 -729 902 -723
rect 904 -729 905 -723
rect 613 -746 617 -740
rect 619 -746 623 -740
rect 358 -767 362 -761
rect 364 -767 368 -761
rect 94 -802 98 -796
rect 100 -802 104 -796
rect -94 -819 -93 -813
rect -91 -819 -90 -813
rect 129 -841 133 -829
rect 135 -841 145 -829
rect 147 -841 150 -829
rect 460 -789 461 -783
rect 463 -789 464 -783
rect 397 -811 400 -805
rect 402 -811 403 -805
rect 407 -811 408 -805
rect 410 -811 411 -805
rect 415 -811 416 -805
rect 418 -811 419 -805
rect 423 -811 424 -805
rect 426 -811 429 -805
rect 539 -807 540 -801
rect 542 -807 543 -801
rect 172 -841 176 -835
rect 178 -841 182 -835
rect -205 -926 -202 -920
rect -200 -926 -185 -920
rect -167 -926 -164 -914
rect -162 -926 -152 -914
rect -150 -926 -147 -914
rect -130 -926 -127 -914
rect -125 -926 -115 -914
rect -113 -926 -110 -914
rect 20 -887 21 -881
rect 23 -887 24 -881
rect 51 -886 55 -874
rect 57 -886 67 -874
rect 69 -886 72 -874
rect 297 -861 301 -849
rect 303 -861 313 -849
rect 315 -861 325 -849
rect 327 -861 328 -849
rect 570 -824 574 -812
rect 576 -824 586 -812
rect 588 -824 591 -812
rect 658 -790 661 -784
rect 663 -790 664 -784
rect 668 -790 669 -784
rect 671 -790 674 -784
rect 698 -790 699 -784
rect 701 -790 702 -784
rect 613 -824 617 -818
rect 619 -824 623 -818
rect 790 -836 793 -830
rect 795 -836 810 -830
rect 828 -836 831 -824
rect 833 -836 843 -824
rect 845 -836 848 -824
rect 865 -836 868 -824
rect 870 -836 880 -824
rect 882 -836 885 -824
rect 901 -836 902 -830
rect 904 -836 905 -830
rect 351 -858 355 -852
rect 357 -858 361 -852
rect 94 -886 98 -880
rect 100 -886 104 -880
rect -94 -926 -93 -920
rect -91 -926 -90 -920
rect 20 -947 21 -941
rect 23 -947 24 -941
rect 51 -964 55 -952
rect 57 -964 67 -952
rect 69 -964 72 -952
rect 136 -930 139 -924
rect 141 -930 142 -924
rect 146 -930 147 -924
rect 149 -930 152 -924
rect 176 -930 177 -924
rect 179 -930 180 -924
rect 297 -947 301 -935
rect 303 -947 313 -935
rect 315 -947 318 -935
rect 540 -912 541 -906
rect 543 -912 544 -906
rect 571 -911 575 -899
rect 577 -911 587 -899
rect 589 -911 592 -899
rect 614 -911 618 -905
rect 620 -911 624 -905
rect 340 -947 344 -941
rect 346 -947 350 -941
rect 790 -943 793 -937
rect 795 -943 810 -937
rect 828 -943 831 -931
rect 833 -943 843 -931
rect 845 -943 848 -931
rect 865 -943 868 -931
rect 870 -943 880 -931
rect 882 -943 885 -931
rect 901 -943 902 -937
rect 904 -943 905 -937
rect 94 -964 98 -958
rect 100 -964 104 -958
rect -205 -1033 -202 -1027
rect -200 -1033 -185 -1027
rect -167 -1033 -164 -1021
rect -162 -1033 -152 -1021
rect -150 -1033 -147 -1021
rect -130 -1033 -127 -1021
rect -125 -1033 -115 -1021
rect -113 -1033 -110 -1021
rect 126 -1003 130 -991
rect 132 -1003 142 -991
rect 144 -1003 147 -991
rect 540 -972 541 -966
rect 543 -972 544 -966
rect 571 -989 575 -977
rect 577 -989 587 -977
rect 589 -989 592 -977
rect 659 -955 662 -949
rect 664 -955 665 -949
rect 669 -955 670 -949
rect 672 -955 675 -949
rect 699 -955 700 -949
rect 702 -955 703 -949
rect 614 -989 618 -983
rect 620 -989 624 -983
rect 169 -1003 173 -997
rect 175 -1003 179 -997
rect -94 -1033 -93 -1027
rect -91 -1033 -90 -1027
rect -205 -1140 -202 -1134
rect -200 -1140 -185 -1134
rect -167 -1140 -164 -1128
rect -162 -1140 -152 -1128
rect -150 -1140 -147 -1128
rect -130 -1140 -127 -1128
rect -125 -1140 -115 -1128
rect -113 -1140 -110 -1128
rect -94 -1140 -93 -1134
rect -91 -1140 -90 -1134
<< pdiffusion >>
rect -205 -240 -202 -216
rect -200 -240 -190 -216
rect -188 -240 -185 -216
rect -167 -228 -164 -216
rect -162 -228 -147 -216
rect -130 -228 -127 -216
rect -125 -228 -110 -216
rect -94 -228 -93 -216
rect -91 -228 -90 -216
rect -205 -347 -202 -323
rect -200 -347 -190 -323
rect -188 -347 -185 -323
rect -167 -335 -164 -323
rect -162 -335 -147 -323
rect -130 -335 -127 -323
rect -125 -335 -110 -323
rect -94 -335 -93 -323
rect -91 -335 -90 -323
rect 54 -361 55 -349
rect 57 -361 60 -349
rect 64 -361 67 -349
rect 69 -361 70 -349
rect 94 -361 98 -349
rect 100 -361 104 -349
rect 20 -379 21 -367
rect 23 -379 24 -367
rect 573 -376 574 -364
rect 576 -376 579 -364
rect 583 -376 586 -364
rect 588 -376 589 -364
rect 613 -376 617 -364
rect 619 -376 623 -364
rect 139 -408 142 -384
rect 144 -408 150 -384
rect 152 -408 155 -384
rect 539 -394 540 -382
rect 542 -394 543 -382
rect -205 -454 -202 -430
rect -200 -454 -190 -430
rect -188 -454 -185 -430
rect -167 -442 -164 -430
rect -162 -442 -147 -430
rect -130 -442 -127 -430
rect -125 -442 -110 -430
rect -94 -442 -93 -430
rect -91 -442 -90 -430
rect 20 -439 21 -427
rect 23 -439 24 -427
rect 54 -439 55 -427
rect 57 -439 60 -427
rect 64 -439 67 -427
rect 69 -439 70 -427
rect 94 -439 98 -427
rect 100 -439 104 -427
rect 179 -422 180 -410
rect 182 -422 183 -410
rect 658 -423 661 -399
rect 663 -423 669 -399
rect 671 -423 674 -399
rect 300 -446 301 -434
rect 303 -446 306 -434
rect 310 -446 313 -434
rect 315 -446 316 -434
rect 340 -446 344 -434
rect 346 -446 350 -434
rect 132 -478 133 -466
rect 135 -478 138 -466
rect 142 -478 145 -466
rect 147 -478 148 -466
rect 172 -478 176 -466
rect 178 -478 182 -466
rect 54 -523 55 -511
rect 57 -523 60 -511
rect 64 -523 67 -511
rect 69 -523 70 -511
rect 94 -523 98 -511
rect 100 -523 104 -511
rect 380 -458 383 -434
rect 385 -458 391 -434
rect 393 -458 396 -434
rect 539 -454 540 -442
rect 542 -454 543 -442
rect 573 -454 574 -442
rect 576 -454 579 -442
rect 583 -454 586 -442
rect 588 -454 589 -442
rect 613 -454 617 -442
rect 619 -454 623 -442
rect 698 -437 699 -425
rect 701 -437 702 -425
rect 420 -472 421 -460
rect 423 -472 424 -460
rect 790 -471 793 -447
rect 795 -471 805 -447
rect 807 -471 810 -447
rect 828 -459 831 -447
rect 833 -459 848 -447
rect 865 -459 868 -447
rect 870 -459 885 -447
rect 901 -459 902 -447
rect 904 -459 905 -447
rect -205 -561 -202 -537
rect -200 -561 -190 -537
rect -188 -561 -185 -537
rect -167 -549 -164 -537
rect -162 -549 -147 -537
rect -130 -549 -127 -537
rect -125 -549 -110 -537
rect -94 -549 -93 -537
rect -91 -549 -90 -537
rect 20 -541 21 -529
rect 23 -541 24 -529
rect 300 -533 301 -521
rect 303 -533 306 -521
rect 310 -533 313 -521
rect 315 -533 318 -521
rect 322 -533 325 -521
rect 327 -533 328 -521
rect 351 -533 355 -521
rect 357 -533 361 -521
rect 136 -570 139 -546
rect 141 -570 147 -546
rect 149 -570 152 -546
rect 20 -601 21 -589
rect 23 -601 24 -589
rect 54 -601 55 -589
rect 57 -601 60 -589
rect 64 -601 67 -589
rect 69 -601 70 -589
rect 94 -601 98 -589
rect 100 -601 104 -589
rect 176 -584 177 -572
rect 179 -584 180 -572
rect 573 -540 574 -528
rect 576 -540 579 -528
rect 583 -540 586 -528
rect 588 -540 589 -528
rect 613 -540 617 -528
rect 619 -540 623 -528
rect 397 -576 400 -552
rect 402 -576 408 -552
rect 410 -576 416 -552
rect 418 -576 421 -552
rect 539 -558 540 -546
rect 542 -558 543 -546
rect 446 -576 447 -564
rect 449 -576 450 -564
rect 658 -587 661 -563
rect 663 -587 669 -563
rect 671 -587 674 -563
rect 790 -578 793 -554
rect 795 -578 805 -554
rect 807 -578 810 -554
rect 828 -566 831 -554
rect 833 -566 848 -554
rect 865 -566 868 -554
rect 870 -566 885 -554
rect 901 -566 902 -554
rect 904 -566 905 -554
rect 300 -628 301 -616
rect 303 -628 306 -616
rect 310 -628 313 -616
rect 315 -628 316 -616
rect 340 -628 344 -616
rect 346 -628 350 -616
rect 539 -618 540 -606
rect 542 -618 543 -606
rect 573 -618 574 -606
rect 576 -618 579 -606
rect 583 -618 586 -606
rect 588 -618 589 -606
rect 613 -618 617 -606
rect 619 -618 623 -606
rect 698 -601 699 -589
rect 701 -601 702 -589
rect 129 -640 130 -628
rect 132 -640 135 -628
rect 139 -640 142 -628
rect 144 -640 145 -628
rect 169 -640 173 -628
rect 175 -640 179 -628
rect -205 -668 -202 -644
rect -200 -668 -190 -644
rect -188 -668 -185 -644
rect -167 -656 -164 -644
rect -162 -656 -147 -644
rect -130 -656 -127 -644
rect -125 -656 -110 -644
rect -94 -656 -93 -644
rect -91 -656 -90 -644
rect 54 -685 55 -673
rect 57 -685 60 -673
rect 64 -685 67 -673
rect 69 -685 70 -673
rect 94 -685 98 -673
rect 100 -685 104 -673
rect 790 -685 793 -661
rect 795 -685 805 -661
rect 807 -685 810 -661
rect 828 -673 831 -661
rect 833 -673 848 -661
rect 865 -673 868 -661
rect 870 -673 885 -661
rect 901 -673 902 -661
rect 904 -673 905 -661
rect 20 -703 21 -691
rect 23 -703 24 -691
rect 139 -732 142 -708
rect 144 -732 150 -708
rect 152 -732 155 -708
rect 300 -717 301 -705
rect 303 -717 306 -705
rect 310 -717 313 -705
rect 315 -717 318 -705
rect 322 -717 325 -705
rect 327 -717 330 -705
rect 334 -717 337 -705
rect 339 -717 340 -705
rect 358 -717 362 -705
rect 364 -717 368 -705
rect 573 -707 574 -695
rect 576 -707 579 -695
rect 583 -707 586 -695
rect 588 -707 589 -695
rect 613 -707 617 -695
rect 619 -707 623 -695
rect -205 -775 -202 -751
rect -200 -775 -190 -751
rect -188 -775 -185 -751
rect -167 -763 -164 -751
rect -162 -763 -147 -751
rect -130 -763 -127 -751
rect -125 -763 -110 -751
rect -94 -763 -93 -751
rect -91 -763 -90 -751
rect 20 -763 21 -751
rect 23 -763 24 -751
rect 54 -763 55 -751
rect 57 -763 60 -751
rect 64 -763 67 -751
rect 69 -763 70 -751
rect 94 -763 98 -751
rect 100 -763 104 -751
rect 179 -746 180 -734
rect 182 -746 183 -734
rect 539 -725 540 -713
rect 542 -725 543 -713
rect 397 -760 400 -736
rect 402 -760 408 -736
rect 410 -760 416 -736
rect 418 -760 424 -736
rect 426 -760 429 -736
rect 658 -754 661 -730
rect 663 -754 669 -730
rect 671 -754 674 -730
rect 132 -802 133 -790
rect 135 -802 138 -790
rect 142 -802 145 -790
rect 147 -802 148 -790
rect 172 -802 176 -790
rect 178 -802 182 -790
rect 54 -847 55 -835
rect 57 -847 60 -835
rect 64 -847 67 -835
rect 69 -847 70 -835
rect 94 -847 98 -835
rect 100 -847 104 -835
rect 300 -815 301 -803
rect 303 -815 306 -803
rect 310 -815 313 -803
rect 315 -815 318 -803
rect 322 -815 325 -803
rect 327 -815 328 -803
rect 351 -815 355 -803
rect 357 -815 361 -803
rect 460 -767 461 -755
rect 463 -767 464 -755
rect 539 -785 540 -773
rect 542 -785 543 -773
rect 573 -785 574 -773
rect 576 -785 579 -773
rect 583 -785 586 -773
rect 588 -785 589 -773
rect 613 -785 617 -773
rect 619 -785 623 -773
rect 698 -768 699 -756
rect 701 -768 702 -756
rect -205 -882 -202 -858
rect -200 -882 -190 -858
rect -188 -882 -185 -858
rect -167 -870 -164 -858
rect -162 -870 -147 -858
rect -130 -870 -127 -858
rect -125 -870 -110 -858
rect -94 -870 -93 -858
rect -91 -870 -90 -858
rect 20 -865 21 -853
rect 23 -865 24 -853
rect 790 -792 793 -768
rect 795 -792 805 -768
rect 807 -792 810 -768
rect 828 -780 831 -768
rect 833 -780 848 -768
rect 865 -780 868 -768
rect 870 -780 885 -768
rect 901 -780 902 -768
rect 904 -780 905 -768
rect 136 -894 139 -870
rect 141 -894 147 -870
rect 149 -894 152 -870
rect 574 -872 575 -860
rect 577 -872 580 -860
rect 584 -872 587 -860
rect 589 -872 590 -860
rect 614 -872 618 -860
rect 620 -872 624 -860
rect 540 -890 541 -878
rect 543 -890 544 -878
rect 20 -925 21 -913
rect 23 -925 24 -913
rect 54 -925 55 -913
rect 57 -925 60 -913
rect 64 -925 67 -913
rect 69 -925 70 -913
rect 94 -925 98 -913
rect 100 -925 104 -913
rect 176 -908 177 -896
rect 179 -908 180 -896
rect 300 -908 301 -896
rect 303 -908 306 -896
rect 310 -908 313 -896
rect 315 -908 316 -896
rect 340 -908 344 -896
rect 346 -908 350 -896
rect 659 -919 662 -895
rect 664 -919 670 -895
rect 672 -919 675 -895
rect 790 -899 793 -875
rect 795 -899 805 -875
rect 807 -899 810 -875
rect 828 -887 831 -875
rect 833 -887 848 -875
rect 865 -887 868 -875
rect 870 -887 885 -875
rect 901 -887 902 -875
rect 904 -887 905 -875
rect 540 -950 541 -938
rect 543 -950 544 -938
rect 574 -950 575 -938
rect 577 -950 580 -938
rect 584 -950 587 -938
rect 589 -950 590 -938
rect 614 -950 618 -938
rect 620 -950 624 -938
rect 699 -933 700 -921
rect 702 -933 703 -921
rect 129 -964 130 -952
rect 132 -964 135 -952
rect 139 -964 142 -952
rect 144 -964 145 -952
rect 169 -964 173 -952
rect 175 -964 179 -952
rect -205 -989 -202 -965
rect -200 -989 -190 -965
rect -188 -989 -185 -965
rect -167 -977 -164 -965
rect -162 -977 -147 -965
rect -130 -977 -127 -965
rect -125 -977 -110 -965
rect -94 -977 -93 -965
rect -91 -977 -90 -965
rect -205 -1096 -202 -1072
rect -200 -1096 -190 -1072
rect -188 -1096 -185 -1072
rect -167 -1084 -164 -1072
rect -162 -1084 -147 -1072
rect -130 -1084 -127 -1072
rect -125 -1084 -110 -1072
rect -94 -1084 -93 -1072
rect -91 -1084 -90 -1072
<< ndcontact >>
rect -209 -284 -205 -278
rect -185 -284 -181 -278
rect -171 -284 -167 -272
rect -147 -284 -143 -272
rect -134 -284 -130 -272
rect -110 -284 -106 -272
rect -98 -284 -94 -278
rect -90 -284 -86 -278
rect -209 -391 -205 -385
rect -185 -391 -181 -385
rect -171 -391 -167 -379
rect -147 -391 -143 -379
rect -134 -391 -130 -379
rect -110 -391 -106 -379
rect -98 -391 -94 -385
rect -90 -391 -86 -385
rect 16 -401 20 -395
rect 24 -401 28 -395
rect 47 -400 51 -388
rect 72 -400 76 -388
rect 90 -400 94 -394
rect 104 -400 108 -394
rect 535 -416 539 -410
rect 543 -416 547 -410
rect 566 -415 570 -403
rect 591 -415 595 -403
rect 609 -415 613 -409
rect 623 -415 627 -409
rect -209 -498 -205 -492
rect -185 -498 -181 -492
rect -171 -498 -167 -486
rect -147 -498 -143 -486
rect -134 -498 -130 -486
rect -110 -498 -106 -486
rect 16 -461 20 -455
rect 24 -461 28 -455
rect 47 -478 51 -466
rect 72 -478 76 -466
rect 135 -444 139 -438
rect 145 -444 149 -438
rect 155 -444 159 -438
rect 175 -444 179 -438
rect 183 -444 187 -438
rect 90 -478 94 -472
rect 104 -478 108 -472
rect -98 -498 -94 -492
rect -90 -498 -86 -492
rect 125 -517 129 -505
rect 150 -517 154 -505
rect 293 -485 297 -473
rect 318 -485 322 -473
rect 336 -485 340 -479
rect 350 -485 354 -479
rect 535 -476 539 -470
rect 543 -476 547 -470
rect 376 -494 380 -488
rect 386 -494 390 -488
rect 396 -494 400 -488
rect 416 -494 420 -488
rect 424 -494 428 -488
rect 566 -493 570 -481
rect 591 -493 595 -481
rect 654 -459 658 -453
rect 664 -459 668 -453
rect 674 -459 678 -453
rect 694 -459 698 -453
rect 702 -459 706 -453
rect 609 -493 613 -487
rect 623 -493 627 -487
rect 168 -517 172 -511
rect 182 -517 186 -511
rect 786 -515 790 -509
rect 810 -515 814 -509
rect 824 -515 828 -503
rect 848 -515 852 -503
rect 861 -515 865 -503
rect 885 -515 889 -503
rect 897 -515 901 -509
rect 905 -515 909 -509
rect -209 -605 -205 -599
rect -185 -605 -181 -599
rect -171 -605 -167 -593
rect -147 -605 -143 -593
rect -134 -605 -130 -593
rect -110 -605 -106 -593
rect 16 -563 20 -557
rect 24 -563 28 -557
rect 47 -562 51 -550
rect 72 -562 76 -550
rect 90 -562 94 -556
rect 104 -562 108 -556
rect -98 -605 -94 -599
rect -90 -605 -86 -599
rect 293 -579 297 -567
rect 328 -579 332 -567
rect 347 -576 351 -570
rect 361 -576 365 -570
rect 16 -623 20 -617
rect 24 -623 28 -617
rect 47 -640 51 -628
rect 72 -640 76 -628
rect 132 -606 136 -600
rect 142 -606 146 -600
rect 152 -606 156 -600
rect 172 -606 176 -600
rect 180 -606 184 -600
rect 535 -580 539 -574
rect 543 -580 547 -574
rect 566 -579 570 -567
rect 591 -579 595 -567
rect 609 -579 613 -573
rect 623 -579 627 -573
rect 442 -598 446 -592
rect 450 -598 454 -592
rect 393 -619 397 -613
rect 403 -619 407 -613
rect 411 -619 415 -613
rect 421 -619 425 -613
rect 90 -640 94 -634
rect 104 -640 108 -634
rect -209 -712 -205 -706
rect -185 -712 -181 -706
rect -171 -712 -167 -700
rect -147 -712 -143 -700
rect -134 -712 -130 -700
rect -110 -712 -106 -700
rect 122 -679 126 -667
rect 147 -679 151 -667
rect 293 -667 297 -655
rect 318 -667 322 -655
rect 535 -640 539 -634
rect 543 -640 547 -634
rect 566 -657 570 -645
rect 591 -657 595 -645
rect 654 -623 658 -617
rect 664 -623 668 -617
rect 674 -623 678 -617
rect 694 -623 698 -617
rect 702 -623 706 -617
rect 786 -622 790 -616
rect 810 -622 814 -616
rect 824 -622 828 -610
rect 848 -622 852 -610
rect 861 -622 865 -610
rect 885 -622 889 -610
rect 897 -622 901 -616
rect 905 -622 909 -616
rect 609 -657 613 -651
rect 623 -657 627 -651
rect 336 -667 340 -661
rect 350 -667 354 -661
rect 165 -679 169 -673
rect 179 -679 183 -673
rect -98 -712 -94 -706
rect -90 -712 -86 -706
rect 16 -725 20 -719
rect 24 -725 28 -719
rect 47 -724 51 -712
rect 72 -724 76 -712
rect 90 -724 94 -718
rect 104 -724 108 -718
rect -209 -819 -205 -813
rect -185 -819 -181 -813
rect -171 -819 -167 -807
rect -147 -819 -143 -807
rect -134 -819 -130 -807
rect -110 -819 -106 -807
rect 16 -785 20 -779
rect 24 -785 28 -779
rect 47 -802 51 -790
rect 72 -802 76 -790
rect 135 -768 139 -762
rect 145 -768 149 -762
rect 155 -768 159 -762
rect 175 -768 179 -762
rect 183 -768 187 -762
rect 293 -770 297 -758
rect 340 -770 344 -758
rect 535 -747 539 -741
rect 543 -747 547 -741
rect 566 -746 570 -734
rect 591 -746 595 -734
rect 786 -729 790 -723
rect 810 -729 814 -723
rect 824 -729 828 -717
rect 848 -729 852 -717
rect 861 -729 865 -717
rect 885 -729 889 -717
rect 897 -729 901 -723
rect 905 -729 909 -723
rect 609 -746 613 -740
rect 623 -746 627 -740
rect 354 -767 358 -761
rect 368 -767 372 -761
rect 90 -802 94 -796
rect 104 -802 108 -796
rect -98 -819 -94 -813
rect -90 -819 -86 -813
rect 125 -841 129 -829
rect 150 -841 154 -829
rect 456 -789 460 -783
rect 464 -789 468 -783
rect 393 -811 397 -805
rect 403 -811 407 -805
rect 411 -811 415 -805
rect 419 -811 423 -805
rect 429 -811 433 -805
rect 535 -807 539 -801
rect 543 -807 547 -801
rect 168 -841 172 -835
rect 182 -841 186 -835
rect -209 -926 -205 -920
rect -185 -926 -181 -920
rect -171 -926 -167 -914
rect -147 -926 -143 -914
rect -134 -926 -130 -914
rect -110 -926 -106 -914
rect 16 -887 20 -881
rect 24 -887 28 -881
rect 47 -886 51 -874
rect 72 -886 76 -874
rect 293 -861 297 -849
rect 328 -861 332 -849
rect 566 -824 570 -812
rect 591 -824 595 -812
rect 654 -790 658 -784
rect 664 -790 668 -784
rect 674 -790 678 -784
rect 694 -790 698 -784
rect 702 -790 706 -784
rect 609 -824 613 -818
rect 623 -824 627 -818
rect 786 -836 790 -830
rect 810 -836 814 -830
rect 824 -836 828 -824
rect 848 -836 852 -824
rect 861 -836 865 -824
rect 885 -836 889 -824
rect 897 -836 901 -830
rect 905 -836 909 -830
rect 347 -858 351 -852
rect 361 -858 365 -852
rect 90 -886 94 -880
rect 104 -886 108 -880
rect -98 -926 -94 -920
rect -90 -926 -86 -920
rect 16 -947 20 -941
rect 24 -947 28 -941
rect 47 -964 51 -952
rect 72 -964 76 -952
rect 132 -930 136 -924
rect 142 -930 146 -924
rect 152 -930 156 -924
rect 172 -930 176 -924
rect 180 -930 184 -924
rect 293 -947 297 -935
rect 318 -947 322 -935
rect 536 -912 540 -906
rect 544 -912 548 -906
rect 567 -911 571 -899
rect 592 -911 596 -899
rect 610 -911 614 -905
rect 624 -911 628 -905
rect 336 -947 340 -941
rect 350 -947 354 -941
rect 786 -943 790 -937
rect 810 -943 814 -937
rect 824 -943 828 -931
rect 848 -943 852 -931
rect 861 -943 865 -931
rect 885 -943 889 -931
rect 897 -943 901 -937
rect 905 -943 909 -937
rect 90 -964 94 -958
rect 104 -964 108 -958
rect -209 -1033 -205 -1027
rect -185 -1033 -181 -1027
rect -171 -1033 -167 -1021
rect -147 -1033 -143 -1021
rect -134 -1033 -130 -1021
rect -110 -1033 -106 -1021
rect 122 -1003 126 -991
rect 147 -1003 151 -991
rect 536 -972 540 -966
rect 544 -972 548 -966
rect 567 -989 571 -977
rect 592 -989 596 -977
rect 655 -955 659 -949
rect 665 -955 669 -949
rect 675 -955 679 -949
rect 695 -955 699 -949
rect 703 -955 707 -949
rect 610 -989 614 -983
rect 624 -989 628 -983
rect 165 -1003 169 -997
rect 179 -1003 183 -997
rect -98 -1033 -94 -1027
rect -90 -1033 -86 -1027
rect -209 -1140 -205 -1134
rect -185 -1140 -181 -1134
rect -171 -1140 -167 -1128
rect -147 -1140 -143 -1128
rect -134 -1140 -130 -1128
rect -110 -1140 -106 -1128
rect -98 -1140 -94 -1134
rect -90 -1140 -86 -1134
<< pdcontact >>
rect -209 -240 -205 -216
rect -185 -240 -181 -216
rect -171 -228 -167 -216
rect -147 -228 -143 -216
rect -134 -228 -130 -216
rect -110 -228 -106 -216
rect -98 -228 -94 -216
rect -90 -228 -86 -216
rect -209 -347 -205 -323
rect -185 -347 -181 -323
rect -171 -335 -167 -323
rect -147 -335 -143 -323
rect -134 -335 -130 -323
rect -110 -335 -106 -323
rect -98 -335 -94 -323
rect -90 -335 -86 -323
rect 50 -361 54 -349
rect 60 -361 64 -349
rect 70 -361 74 -349
rect 90 -361 94 -349
rect 104 -361 108 -349
rect 16 -379 20 -367
rect 24 -379 28 -367
rect 569 -376 573 -364
rect 579 -376 583 -364
rect 589 -376 593 -364
rect 609 -376 613 -364
rect 623 -376 627 -364
rect 135 -408 139 -384
rect 155 -408 159 -384
rect 535 -394 539 -382
rect 543 -394 547 -382
rect -209 -454 -205 -430
rect -185 -454 -181 -430
rect -171 -442 -167 -430
rect -147 -442 -143 -430
rect -134 -442 -130 -430
rect -110 -442 -106 -430
rect -98 -442 -94 -430
rect -90 -442 -86 -430
rect 16 -439 20 -427
rect 24 -439 28 -427
rect 50 -439 54 -427
rect 60 -439 64 -427
rect 70 -439 74 -427
rect 90 -439 94 -427
rect 104 -439 108 -427
rect 175 -422 179 -410
rect 183 -422 187 -410
rect 654 -423 658 -399
rect 674 -423 678 -399
rect 296 -446 300 -434
rect 306 -446 310 -434
rect 316 -446 320 -434
rect 336 -446 340 -434
rect 350 -446 354 -434
rect 128 -478 132 -466
rect 138 -478 142 -466
rect 148 -478 152 -466
rect 168 -478 172 -466
rect 182 -478 186 -466
rect 50 -523 54 -511
rect 60 -523 64 -511
rect 70 -523 74 -511
rect 90 -523 94 -511
rect 104 -523 108 -511
rect 376 -458 380 -434
rect 396 -458 400 -434
rect 535 -454 539 -442
rect 543 -454 547 -442
rect 569 -454 573 -442
rect 579 -454 583 -442
rect 589 -454 593 -442
rect 609 -454 613 -442
rect 623 -454 627 -442
rect 694 -437 698 -425
rect 702 -437 706 -425
rect 416 -472 420 -460
rect 424 -472 428 -460
rect 786 -471 790 -447
rect 810 -471 814 -447
rect 824 -459 828 -447
rect 848 -459 852 -447
rect 861 -459 865 -447
rect 885 -459 889 -447
rect 897 -459 901 -447
rect 905 -459 909 -447
rect -209 -561 -205 -537
rect -185 -561 -181 -537
rect -171 -549 -167 -537
rect -147 -549 -143 -537
rect -134 -549 -130 -537
rect -110 -549 -106 -537
rect -98 -549 -94 -537
rect -90 -549 -86 -537
rect 16 -541 20 -529
rect 24 -541 28 -529
rect 296 -533 300 -521
rect 306 -533 310 -521
rect 318 -533 322 -521
rect 328 -533 332 -521
rect 347 -533 351 -521
rect 361 -533 365 -521
rect 132 -570 136 -546
rect 152 -570 156 -546
rect 16 -601 20 -589
rect 24 -601 28 -589
rect 50 -601 54 -589
rect 60 -601 64 -589
rect 70 -601 74 -589
rect 90 -601 94 -589
rect 104 -601 108 -589
rect 172 -584 176 -572
rect 180 -584 184 -572
rect 569 -540 573 -528
rect 579 -540 583 -528
rect 589 -540 593 -528
rect 609 -540 613 -528
rect 623 -540 627 -528
rect 393 -576 397 -552
rect 421 -576 425 -552
rect 535 -558 539 -546
rect 543 -558 547 -546
rect 442 -576 446 -564
rect 450 -576 454 -564
rect 654 -587 658 -563
rect 674 -587 678 -563
rect 786 -578 790 -554
rect 810 -578 814 -554
rect 824 -566 828 -554
rect 848 -566 852 -554
rect 861 -566 865 -554
rect 885 -566 889 -554
rect 897 -566 901 -554
rect 905 -566 909 -554
rect 296 -628 300 -616
rect 306 -628 310 -616
rect 316 -628 320 -616
rect 336 -628 340 -616
rect 350 -628 354 -616
rect 535 -618 539 -606
rect 543 -618 547 -606
rect 569 -618 573 -606
rect 579 -618 583 -606
rect 589 -618 593 -606
rect 609 -618 613 -606
rect 623 -618 627 -606
rect 694 -601 698 -589
rect 702 -601 706 -589
rect 125 -640 129 -628
rect 135 -640 139 -628
rect 145 -640 149 -628
rect 165 -640 169 -628
rect 179 -640 183 -628
rect -209 -668 -205 -644
rect -185 -668 -181 -644
rect -171 -656 -167 -644
rect -147 -656 -143 -644
rect -134 -656 -130 -644
rect -110 -656 -106 -644
rect -98 -656 -94 -644
rect -90 -656 -86 -644
rect 50 -685 54 -673
rect 60 -685 64 -673
rect 70 -685 74 -673
rect 90 -685 94 -673
rect 104 -685 108 -673
rect 786 -685 790 -661
rect 810 -685 814 -661
rect 824 -673 828 -661
rect 848 -673 852 -661
rect 861 -673 865 -661
rect 885 -673 889 -661
rect 897 -673 901 -661
rect 905 -673 909 -661
rect 16 -703 20 -691
rect 24 -703 28 -691
rect 135 -732 139 -708
rect 155 -732 159 -708
rect 296 -717 300 -705
rect 306 -717 310 -705
rect 318 -717 322 -705
rect 330 -717 334 -705
rect 340 -717 344 -705
rect 354 -717 358 -705
rect 368 -717 372 -705
rect 569 -707 573 -695
rect 579 -707 583 -695
rect 589 -707 593 -695
rect 609 -707 613 -695
rect 623 -707 627 -695
rect -209 -775 -205 -751
rect -185 -775 -181 -751
rect -171 -763 -167 -751
rect -147 -763 -143 -751
rect -134 -763 -130 -751
rect -110 -763 -106 -751
rect -98 -763 -94 -751
rect -90 -763 -86 -751
rect 16 -763 20 -751
rect 24 -763 28 -751
rect 50 -763 54 -751
rect 60 -763 64 -751
rect 70 -763 74 -751
rect 90 -763 94 -751
rect 104 -763 108 -751
rect 175 -746 179 -734
rect 183 -746 187 -734
rect 535 -725 539 -713
rect 543 -725 547 -713
rect 393 -760 397 -736
rect 429 -760 433 -736
rect 654 -754 658 -730
rect 674 -754 678 -730
rect 128 -802 132 -790
rect 138 -802 142 -790
rect 148 -802 152 -790
rect 168 -802 172 -790
rect 182 -802 186 -790
rect 50 -847 54 -835
rect 60 -847 64 -835
rect 70 -847 74 -835
rect 90 -847 94 -835
rect 104 -847 108 -835
rect 296 -815 300 -803
rect 306 -815 310 -803
rect 318 -815 322 -803
rect 328 -815 332 -803
rect 347 -815 351 -803
rect 361 -815 365 -803
rect 456 -767 460 -755
rect 464 -767 468 -755
rect 535 -785 539 -773
rect 543 -785 547 -773
rect 569 -785 573 -773
rect 579 -785 583 -773
rect 589 -785 593 -773
rect 609 -785 613 -773
rect 623 -785 627 -773
rect 694 -768 698 -756
rect 702 -768 706 -756
rect -209 -882 -205 -858
rect -185 -882 -181 -858
rect -171 -870 -167 -858
rect -147 -870 -143 -858
rect -134 -870 -130 -858
rect -110 -870 -106 -858
rect -98 -870 -94 -858
rect -90 -870 -86 -858
rect 16 -865 20 -853
rect 24 -865 28 -853
rect 786 -792 790 -768
rect 810 -792 814 -768
rect 824 -780 828 -768
rect 848 -780 852 -768
rect 861 -780 865 -768
rect 885 -780 889 -768
rect 897 -780 901 -768
rect 905 -780 909 -768
rect 132 -894 136 -870
rect 152 -894 156 -870
rect 570 -872 574 -860
rect 580 -872 584 -860
rect 590 -872 594 -860
rect 610 -872 614 -860
rect 624 -872 628 -860
rect 536 -890 540 -878
rect 544 -890 548 -878
rect 16 -925 20 -913
rect 24 -925 28 -913
rect 50 -925 54 -913
rect 60 -925 64 -913
rect 70 -925 74 -913
rect 90 -925 94 -913
rect 104 -925 108 -913
rect 172 -908 176 -896
rect 180 -908 184 -896
rect 296 -908 300 -896
rect 306 -908 310 -896
rect 316 -908 320 -896
rect 336 -908 340 -896
rect 350 -908 354 -896
rect 655 -919 659 -895
rect 675 -919 679 -895
rect 786 -899 790 -875
rect 810 -899 814 -875
rect 824 -887 828 -875
rect 848 -887 852 -875
rect 861 -887 865 -875
rect 885 -887 889 -875
rect 897 -887 901 -875
rect 905 -887 909 -875
rect 536 -950 540 -938
rect 544 -950 548 -938
rect 570 -950 574 -938
rect 580 -950 584 -938
rect 590 -950 594 -938
rect 610 -950 614 -938
rect 624 -950 628 -938
rect 695 -933 699 -921
rect 703 -933 707 -921
rect 125 -964 129 -952
rect 135 -964 139 -952
rect 145 -964 149 -952
rect 165 -964 169 -952
rect 179 -964 183 -952
rect -209 -989 -205 -965
rect -185 -989 -181 -965
rect -171 -977 -167 -965
rect -147 -977 -143 -965
rect -134 -977 -130 -965
rect -110 -977 -106 -965
rect -98 -977 -94 -965
rect -90 -977 -86 -965
rect -209 -1096 -205 -1072
rect -185 -1096 -181 -1072
rect -171 -1084 -167 -1072
rect -147 -1084 -143 -1072
rect -134 -1084 -130 -1072
rect -110 -1084 -106 -1072
rect -98 -1084 -94 -1072
rect -90 -1084 -86 -1072
<< polysilicon >>
rect -202 -216 -200 -213
rect -190 -216 -188 -213
rect -164 -216 -162 -213
rect -127 -216 -125 -213
rect -93 -216 -91 -213
rect -202 -278 -200 -240
rect -190 -258 -188 -240
rect -164 -272 -162 -240
rect -152 -272 -150 -262
rect -127 -272 -125 -240
rect -115 -272 -113 -254
rect -93 -278 -91 -228
rect -202 -287 -200 -284
rect -164 -287 -162 -284
rect -152 -287 -150 -284
rect -127 -287 -125 -284
rect -115 -287 -113 -284
rect -93 -287 -91 -284
rect -202 -323 -200 -320
rect -190 -323 -188 -320
rect -164 -323 -162 -320
rect -127 -323 -125 -320
rect -93 -323 -91 -320
rect -202 -385 -200 -347
rect -190 -365 -188 -347
rect -164 -379 -162 -347
rect -152 -379 -150 -369
rect -127 -379 -125 -347
rect -115 -379 -113 -361
rect -93 -385 -91 -335
rect 55 -349 57 -346
rect 67 -349 69 -346
rect 98 -349 100 -346
rect 21 -367 23 -364
rect -202 -394 -200 -391
rect -164 -394 -162 -391
rect -152 -394 -150 -391
rect -127 -394 -125 -391
rect -115 -394 -113 -391
rect -93 -394 -91 -391
rect 21 -395 23 -379
rect 55 -388 57 -361
rect 67 -388 69 -361
rect 98 -394 100 -361
rect 574 -364 576 -361
rect 586 -364 588 -361
rect 617 -364 619 -361
rect 142 -384 144 -381
rect 150 -384 152 -381
rect 540 -382 542 -379
rect 21 -404 23 -401
rect 55 -403 57 -400
rect 67 -403 69 -400
rect 98 -403 100 -400
rect 142 -417 144 -408
rect 21 -427 23 -424
rect 55 -427 57 -424
rect 67 -427 69 -424
rect 98 -427 100 -424
rect -202 -430 -200 -427
rect -190 -430 -188 -427
rect -164 -430 -162 -427
rect -127 -430 -125 -427
rect -93 -430 -91 -427
rect 142 -438 144 -421
rect 150 -424 152 -408
rect 180 -410 182 -407
rect 540 -410 542 -394
rect 574 -403 576 -376
rect 586 -403 588 -376
rect 617 -409 619 -376
rect 661 -399 663 -396
rect 669 -399 671 -396
rect 540 -419 542 -416
rect 574 -418 576 -415
rect 586 -418 588 -415
rect 617 -418 619 -415
rect 150 -438 152 -428
rect 180 -438 182 -422
rect 301 -434 303 -431
rect 313 -434 315 -431
rect 344 -434 346 -431
rect 383 -434 385 -431
rect 391 -434 393 -431
rect 661 -432 663 -423
rect -202 -492 -200 -454
rect -190 -472 -188 -454
rect -164 -486 -162 -454
rect -152 -486 -150 -476
rect -127 -486 -125 -454
rect -115 -486 -113 -468
rect -93 -492 -91 -442
rect 21 -455 23 -439
rect 21 -464 23 -461
rect 55 -466 57 -439
rect 67 -466 69 -439
rect 98 -472 100 -439
rect 142 -447 144 -444
rect 150 -447 152 -444
rect 180 -448 182 -444
rect 133 -466 135 -463
rect 145 -466 147 -463
rect 176 -466 178 -463
rect 301 -473 303 -446
rect 313 -473 315 -446
rect 55 -481 57 -478
rect 67 -481 69 -478
rect 98 -481 100 -478
rect -202 -501 -200 -498
rect -164 -501 -162 -498
rect -152 -501 -150 -498
rect -127 -501 -125 -498
rect -115 -501 -113 -498
rect -93 -501 -91 -498
rect 133 -505 135 -478
rect 145 -505 147 -478
rect 55 -511 57 -508
rect 67 -511 69 -508
rect 98 -511 100 -508
rect 176 -511 178 -478
rect 344 -479 346 -446
rect 540 -442 542 -439
rect 574 -442 576 -439
rect 586 -442 588 -439
rect 617 -442 619 -439
rect 661 -453 663 -436
rect 669 -439 671 -423
rect 699 -425 701 -422
rect 669 -453 671 -443
rect 699 -453 701 -437
rect 793 -447 795 -444
rect 805 -447 807 -444
rect 831 -447 833 -444
rect 868 -447 870 -444
rect 902 -447 904 -444
rect 383 -467 385 -458
rect 301 -488 303 -485
rect 313 -488 315 -485
rect 344 -488 346 -485
rect 383 -488 385 -471
rect 391 -474 393 -458
rect 421 -460 423 -457
rect 540 -470 542 -454
rect 391 -488 393 -478
rect 421 -488 423 -472
rect 540 -479 542 -476
rect 574 -481 576 -454
rect 586 -481 588 -454
rect 617 -487 619 -454
rect 661 -462 663 -459
rect 669 -462 671 -459
rect 699 -463 701 -459
rect 383 -497 385 -494
rect 391 -497 393 -494
rect 421 -498 423 -494
rect 574 -496 576 -493
rect 586 -496 588 -493
rect 617 -496 619 -493
rect 793 -509 795 -471
rect 805 -489 807 -471
rect 831 -503 833 -471
rect 843 -503 845 -493
rect 868 -503 870 -471
rect 880 -503 882 -485
rect 902 -509 904 -459
rect 133 -520 135 -517
rect 145 -520 147 -517
rect 176 -520 178 -517
rect 793 -518 795 -515
rect 831 -518 833 -515
rect 843 -518 845 -515
rect 868 -518 870 -515
rect 880 -518 882 -515
rect 902 -518 904 -515
rect 301 -521 303 -518
rect 313 -521 315 -518
rect 325 -521 327 -518
rect 355 -521 357 -518
rect 21 -529 23 -526
rect -202 -537 -200 -534
rect -190 -537 -188 -534
rect -164 -537 -162 -534
rect -127 -537 -125 -534
rect -93 -537 -91 -534
rect -202 -599 -200 -561
rect -190 -579 -188 -561
rect -164 -593 -162 -561
rect -152 -593 -150 -583
rect -127 -593 -125 -561
rect -115 -593 -113 -575
rect -93 -599 -91 -549
rect 21 -557 23 -541
rect 55 -550 57 -523
rect 67 -550 69 -523
rect 98 -556 100 -523
rect 574 -528 576 -525
rect 586 -528 588 -525
rect 617 -528 619 -525
rect 139 -546 141 -543
rect 147 -546 149 -543
rect 21 -566 23 -563
rect 55 -565 57 -562
rect 67 -565 69 -562
rect 98 -565 100 -562
rect 301 -567 303 -533
rect 313 -567 315 -533
rect 325 -567 327 -533
rect 139 -579 141 -570
rect 21 -589 23 -586
rect 55 -589 57 -586
rect 67 -589 69 -586
rect 98 -589 100 -586
rect 139 -600 141 -583
rect 147 -586 149 -570
rect 177 -572 179 -569
rect 355 -570 357 -533
rect 540 -546 542 -543
rect 400 -552 402 -549
rect 408 -552 410 -549
rect 416 -552 418 -549
rect 447 -564 449 -561
rect 540 -574 542 -558
rect 574 -567 576 -540
rect 586 -567 588 -540
rect 355 -579 357 -576
rect 301 -582 303 -579
rect 313 -582 315 -579
rect 325 -582 327 -579
rect 147 -600 149 -590
rect 177 -600 179 -584
rect 400 -585 402 -576
rect -202 -608 -200 -605
rect -164 -608 -162 -605
rect -152 -608 -150 -605
rect -127 -608 -125 -605
rect -115 -608 -113 -605
rect -93 -608 -91 -605
rect 21 -617 23 -601
rect 21 -626 23 -623
rect 55 -628 57 -601
rect 67 -628 69 -601
rect 98 -634 100 -601
rect 139 -609 141 -606
rect 147 -609 149 -606
rect 177 -610 179 -606
rect 400 -613 402 -589
rect 408 -592 410 -576
rect 408 -613 410 -596
rect 416 -599 418 -576
rect 447 -592 449 -576
rect 617 -573 619 -540
rect 793 -554 795 -551
rect 805 -554 807 -551
rect 831 -554 833 -551
rect 868 -554 870 -551
rect 902 -554 904 -551
rect 661 -563 663 -560
rect 669 -563 671 -560
rect 540 -583 542 -580
rect 574 -582 576 -579
rect 586 -582 588 -579
rect 617 -582 619 -579
rect 661 -596 663 -587
rect 447 -601 449 -598
rect 416 -613 418 -603
rect 540 -606 542 -603
rect 574 -606 576 -603
rect 586 -606 588 -603
rect 617 -606 619 -603
rect 301 -616 303 -613
rect 313 -616 315 -613
rect 344 -616 346 -613
rect 130 -628 132 -625
rect 142 -628 144 -625
rect 173 -628 175 -625
rect 661 -617 663 -600
rect 669 -603 671 -587
rect 699 -589 701 -586
rect 669 -617 671 -607
rect 699 -617 701 -601
rect 793 -616 795 -578
rect 805 -596 807 -578
rect 831 -610 833 -578
rect 843 -610 845 -600
rect 868 -610 870 -578
rect 880 -610 882 -592
rect 400 -622 402 -619
rect 408 -622 410 -619
rect 416 -622 418 -619
rect -202 -644 -200 -641
rect -190 -644 -188 -641
rect -164 -644 -162 -641
rect -127 -644 -125 -641
rect -93 -644 -91 -641
rect 55 -643 57 -640
rect 67 -643 69 -640
rect 98 -643 100 -640
rect -202 -706 -200 -668
rect -190 -686 -188 -668
rect -164 -700 -162 -668
rect -152 -700 -150 -690
rect -127 -700 -125 -668
rect -115 -700 -113 -682
rect -93 -706 -91 -656
rect 130 -667 132 -640
rect 142 -667 144 -640
rect 55 -673 57 -670
rect 67 -673 69 -670
rect 98 -673 100 -670
rect 173 -673 175 -640
rect 301 -655 303 -628
rect 313 -655 315 -628
rect 344 -661 346 -628
rect 540 -634 542 -618
rect 540 -643 542 -640
rect 574 -645 576 -618
rect 586 -645 588 -618
rect 617 -651 619 -618
rect 902 -616 904 -566
rect 661 -626 663 -623
rect 669 -626 671 -623
rect 699 -627 701 -623
rect 793 -625 795 -622
rect 831 -625 833 -622
rect 843 -625 845 -622
rect 868 -625 870 -622
rect 880 -625 882 -622
rect 902 -625 904 -622
rect 574 -660 576 -657
rect 586 -660 588 -657
rect 617 -660 619 -657
rect 793 -661 795 -658
rect 805 -661 807 -658
rect 831 -661 833 -658
rect 868 -661 870 -658
rect 902 -661 904 -658
rect 301 -670 303 -667
rect 313 -670 315 -667
rect 344 -670 346 -667
rect 130 -682 132 -679
rect 142 -682 144 -679
rect 173 -682 175 -679
rect 21 -691 23 -688
rect -202 -715 -200 -712
rect -164 -715 -162 -712
rect -152 -715 -150 -712
rect -127 -715 -125 -712
rect -115 -715 -113 -712
rect -93 -715 -91 -712
rect 21 -719 23 -703
rect 55 -712 57 -685
rect 67 -712 69 -685
rect 98 -718 100 -685
rect 574 -695 576 -692
rect 586 -695 588 -692
rect 617 -695 619 -692
rect 301 -705 303 -702
rect 313 -705 315 -702
rect 325 -705 327 -702
rect 337 -705 339 -702
rect 362 -705 364 -702
rect 142 -708 144 -705
rect 150 -708 152 -705
rect 21 -728 23 -725
rect 55 -727 57 -724
rect 67 -727 69 -724
rect 98 -727 100 -724
rect 540 -713 542 -710
rect 142 -741 144 -732
rect -202 -751 -200 -748
rect -190 -751 -188 -748
rect -164 -751 -162 -748
rect -127 -751 -125 -748
rect -93 -751 -91 -748
rect 21 -751 23 -748
rect 55 -751 57 -748
rect 67 -751 69 -748
rect 98 -751 100 -748
rect 142 -762 144 -745
rect 150 -748 152 -732
rect 180 -734 182 -731
rect 150 -762 152 -752
rect 180 -762 182 -746
rect 301 -758 303 -717
rect 313 -758 315 -717
rect 325 -758 327 -717
rect 337 -758 339 -717
rect -202 -813 -200 -775
rect -190 -793 -188 -775
rect -164 -807 -162 -775
rect -152 -807 -150 -797
rect -127 -807 -125 -775
rect -115 -807 -113 -789
rect -93 -813 -91 -763
rect 21 -779 23 -763
rect 21 -788 23 -785
rect 55 -790 57 -763
rect 67 -790 69 -763
rect 98 -796 100 -763
rect 142 -771 144 -768
rect 150 -771 152 -768
rect 180 -772 182 -768
rect 362 -761 364 -717
rect 400 -736 402 -733
rect 408 -736 410 -733
rect 416 -736 418 -733
rect 424 -736 426 -733
rect 540 -741 542 -725
rect 574 -734 576 -707
rect 586 -734 588 -707
rect 617 -740 619 -707
rect 793 -723 795 -685
rect 805 -703 807 -685
rect 831 -717 833 -685
rect 843 -717 845 -707
rect 868 -717 870 -685
rect 880 -717 882 -699
rect 661 -730 663 -727
rect 669 -730 671 -727
rect 902 -723 904 -673
rect 540 -750 542 -747
rect 574 -749 576 -746
rect 586 -749 588 -746
rect 617 -749 619 -746
rect 461 -755 463 -752
rect 793 -732 795 -729
rect 831 -732 833 -729
rect 843 -732 845 -729
rect 868 -732 870 -729
rect 880 -732 882 -729
rect 902 -732 904 -729
rect 362 -770 364 -767
rect 400 -769 402 -760
rect 301 -773 303 -770
rect 313 -773 315 -770
rect 325 -773 327 -770
rect 337 -773 339 -770
rect 133 -790 135 -787
rect 145 -790 147 -787
rect 176 -790 178 -787
rect 55 -805 57 -802
rect 67 -805 69 -802
rect 98 -805 100 -802
rect -202 -822 -200 -819
rect -164 -822 -162 -819
rect -152 -822 -150 -819
rect -127 -822 -125 -819
rect -115 -822 -113 -819
rect -93 -822 -91 -819
rect 133 -829 135 -802
rect 145 -829 147 -802
rect 55 -835 57 -832
rect 67 -835 69 -832
rect 98 -835 100 -832
rect 176 -835 178 -802
rect 301 -803 303 -800
rect 313 -803 315 -800
rect 325 -803 327 -800
rect 355 -803 357 -800
rect 400 -805 402 -773
rect 408 -776 410 -760
rect 408 -805 410 -780
rect 416 -783 418 -760
rect 416 -805 418 -787
rect 424 -790 426 -760
rect 661 -763 663 -754
rect 461 -783 463 -767
rect 540 -773 542 -770
rect 574 -773 576 -770
rect 586 -773 588 -770
rect 617 -773 619 -770
rect 661 -784 663 -767
rect 669 -770 671 -754
rect 699 -756 701 -753
rect 793 -768 795 -765
rect 805 -768 807 -765
rect 831 -768 833 -765
rect 868 -768 870 -765
rect 902 -768 904 -765
rect 669 -784 671 -774
rect 699 -784 701 -768
rect 461 -793 463 -789
rect 424 -805 426 -794
rect 540 -801 542 -785
rect 540 -810 542 -807
rect 400 -814 402 -811
rect 408 -814 410 -811
rect 416 -814 418 -811
rect 424 -814 426 -811
rect 574 -812 576 -785
rect 586 -812 588 -785
rect 133 -844 135 -841
rect 145 -844 147 -841
rect 176 -844 178 -841
rect 21 -853 23 -850
rect -202 -858 -200 -855
rect -190 -858 -188 -855
rect -164 -858 -162 -855
rect -127 -858 -125 -855
rect -93 -858 -91 -855
rect -202 -920 -200 -882
rect -190 -900 -188 -882
rect -164 -914 -162 -882
rect -152 -914 -150 -904
rect -127 -914 -125 -882
rect -115 -914 -113 -896
rect -93 -920 -91 -870
rect 21 -881 23 -865
rect 55 -874 57 -847
rect 67 -874 69 -847
rect 98 -880 100 -847
rect 301 -849 303 -815
rect 313 -849 315 -815
rect 325 -849 327 -815
rect 355 -852 357 -815
rect 617 -818 619 -785
rect 661 -793 663 -790
rect 669 -793 671 -790
rect 699 -794 701 -790
rect 574 -827 576 -824
rect 586 -827 588 -824
rect 617 -827 619 -824
rect 793 -830 795 -792
rect 805 -810 807 -792
rect 831 -824 833 -792
rect 843 -824 845 -814
rect 868 -824 870 -792
rect 880 -824 882 -806
rect 902 -830 904 -780
rect 793 -839 795 -836
rect 831 -839 833 -836
rect 843 -839 845 -836
rect 868 -839 870 -836
rect 880 -839 882 -836
rect 902 -839 904 -836
rect 355 -861 357 -858
rect 575 -860 577 -857
rect 587 -860 589 -857
rect 618 -860 620 -857
rect 301 -864 303 -861
rect 313 -864 315 -861
rect 325 -864 327 -861
rect 139 -870 141 -867
rect 147 -870 149 -867
rect 21 -890 23 -887
rect 55 -889 57 -886
rect 67 -889 69 -886
rect 98 -889 100 -886
rect 541 -878 543 -875
rect 139 -903 141 -894
rect 21 -913 23 -910
rect 55 -913 57 -910
rect 67 -913 69 -910
rect 98 -913 100 -910
rect 139 -924 141 -907
rect 147 -910 149 -894
rect 177 -896 179 -893
rect 301 -896 303 -893
rect 313 -896 315 -893
rect 344 -896 346 -893
rect 541 -906 543 -890
rect 575 -899 577 -872
rect 587 -899 589 -872
rect 147 -924 149 -914
rect 177 -924 179 -908
rect -202 -929 -200 -926
rect -164 -929 -162 -926
rect -152 -929 -150 -926
rect -127 -929 -125 -926
rect -115 -929 -113 -926
rect -93 -929 -91 -926
rect 21 -941 23 -925
rect 21 -950 23 -947
rect 55 -952 57 -925
rect 67 -952 69 -925
rect -202 -965 -200 -962
rect -190 -965 -188 -962
rect -164 -965 -162 -962
rect -127 -965 -125 -962
rect -93 -965 -91 -962
rect 98 -958 100 -925
rect 139 -933 141 -930
rect 147 -933 149 -930
rect 177 -934 179 -930
rect 301 -935 303 -908
rect 313 -935 315 -908
rect 344 -941 346 -908
rect 618 -905 620 -872
rect 793 -875 795 -872
rect 805 -875 807 -872
rect 831 -875 833 -872
rect 868 -875 870 -872
rect 902 -875 904 -872
rect 662 -895 664 -892
rect 670 -895 672 -892
rect 541 -915 543 -912
rect 575 -914 577 -911
rect 587 -914 589 -911
rect 618 -914 620 -911
rect 662 -928 664 -919
rect 541 -938 543 -935
rect 575 -938 577 -935
rect 587 -938 589 -935
rect 618 -938 620 -935
rect 130 -952 132 -949
rect 142 -952 144 -949
rect 173 -952 175 -949
rect 301 -950 303 -947
rect 313 -950 315 -947
rect 344 -950 346 -947
rect 662 -949 664 -932
rect 670 -935 672 -919
rect 700 -921 702 -918
rect 670 -949 672 -939
rect 700 -949 702 -933
rect 793 -937 795 -899
rect 805 -917 807 -899
rect 831 -931 833 -899
rect 843 -931 845 -921
rect 868 -931 870 -899
rect 880 -931 882 -913
rect 902 -937 904 -887
rect 793 -946 795 -943
rect 831 -946 833 -943
rect 843 -946 845 -943
rect 868 -946 870 -943
rect 880 -946 882 -943
rect 902 -946 904 -943
rect 55 -967 57 -964
rect 67 -967 69 -964
rect 98 -967 100 -964
rect -202 -1027 -200 -989
rect -190 -1007 -188 -989
rect -164 -1021 -162 -989
rect -152 -1021 -150 -1011
rect -127 -1021 -125 -989
rect -115 -1021 -113 -1003
rect -93 -1027 -91 -977
rect 130 -991 132 -964
rect 142 -991 144 -964
rect 173 -997 175 -964
rect 541 -966 543 -950
rect 541 -975 543 -972
rect 575 -977 577 -950
rect 587 -977 589 -950
rect 618 -983 620 -950
rect 662 -958 664 -955
rect 670 -958 672 -955
rect 700 -959 702 -955
rect 575 -992 577 -989
rect 587 -992 589 -989
rect 618 -992 620 -989
rect 130 -1006 132 -1003
rect 142 -1006 144 -1003
rect 173 -1006 175 -1003
rect -202 -1036 -200 -1033
rect -164 -1036 -162 -1033
rect -152 -1036 -150 -1033
rect -127 -1036 -125 -1033
rect -115 -1036 -113 -1033
rect -93 -1036 -91 -1033
rect -202 -1072 -200 -1069
rect -190 -1072 -188 -1069
rect -164 -1072 -162 -1069
rect -127 -1072 -125 -1069
rect -93 -1072 -91 -1069
rect -202 -1134 -200 -1096
rect -190 -1114 -188 -1096
rect -164 -1128 -162 -1096
rect -152 -1128 -150 -1118
rect -127 -1128 -125 -1096
rect -115 -1128 -113 -1110
rect -93 -1134 -91 -1084
rect -202 -1143 -200 -1140
rect -164 -1143 -162 -1140
rect -152 -1143 -150 -1140
rect -127 -1143 -125 -1140
rect -115 -1143 -113 -1140
rect -93 -1143 -91 -1140
<< polycontact >>
rect -206 -251 -202 -247
rect -194 -258 -190 -254
rect -168 -251 -164 -247
rect -131 -251 -127 -247
rect -156 -266 -152 -262
rect -97 -251 -93 -247
rect -119 -258 -115 -254
rect -206 -358 -202 -354
rect -194 -365 -190 -361
rect -168 -358 -164 -354
rect -131 -358 -127 -354
rect -156 -373 -152 -369
rect -97 -358 -93 -354
rect -119 -365 -115 -361
rect 51 -376 55 -372
rect 17 -392 21 -388
rect 63 -379 67 -375
rect 94 -372 98 -368
rect 570 -391 574 -387
rect 536 -407 540 -403
rect 140 -421 144 -417
rect 582 -394 586 -390
rect 613 -387 617 -383
rect 148 -428 152 -424
rect 176 -435 180 -431
rect -206 -465 -202 -461
rect -194 -472 -190 -468
rect -168 -465 -164 -461
rect -131 -465 -127 -461
rect -156 -480 -152 -476
rect -97 -465 -93 -461
rect -119 -472 -115 -468
rect 17 -452 21 -448
rect 51 -456 55 -452
rect 63 -463 67 -459
rect 94 -452 98 -448
rect 297 -463 301 -459
rect 309 -470 313 -466
rect 340 -459 344 -455
rect 129 -495 133 -491
rect 141 -502 145 -498
rect 172 -491 176 -487
rect 659 -436 663 -432
rect 667 -443 671 -439
rect 695 -450 699 -446
rect 381 -471 385 -467
rect 536 -467 540 -463
rect 389 -478 393 -474
rect 417 -485 421 -481
rect 570 -471 574 -467
rect 582 -478 586 -474
rect 613 -467 617 -463
rect 789 -482 793 -478
rect 801 -489 805 -485
rect 827 -482 831 -478
rect 864 -482 868 -478
rect 839 -497 843 -493
rect 898 -482 902 -478
rect 876 -489 880 -485
rect 51 -538 55 -534
rect -206 -572 -202 -568
rect -194 -579 -190 -575
rect -168 -572 -164 -568
rect -131 -572 -127 -568
rect -156 -587 -152 -583
rect -97 -572 -93 -568
rect -119 -579 -115 -575
rect 17 -554 21 -550
rect 63 -541 67 -537
rect 94 -534 98 -530
rect 297 -550 301 -546
rect 309 -557 313 -553
rect 321 -564 325 -560
rect 351 -546 355 -542
rect 137 -583 141 -579
rect 570 -555 574 -551
rect 536 -571 540 -567
rect 582 -558 586 -554
rect 613 -551 617 -547
rect 145 -590 149 -586
rect 173 -597 177 -593
rect 398 -589 402 -585
rect 17 -614 21 -610
rect 51 -618 55 -614
rect 63 -625 67 -621
rect 94 -614 98 -610
rect 406 -596 410 -592
rect 443 -589 447 -585
rect 414 -603 418 -599
rect 659 -600 663 -596
rect 789 -589 793 -585
rect 667 -607 671 -603
rect 695 -614 699 -610
rect 801 -596 805 -592
rect 827 -589 831 -585
rect 864 -589 868 -585
rect 839 -604 843 -600
rect 898 -589 902 -585
rect 876 -596 880 -592
rect -206 -679 -202 -675
rect -194 -686 -190 -682
rect -168 -679 -164 -675
rect -131 -679 -127 -675
rect -156 -694 -152 -690
rect -97 -679 -93 -675
rect -119 -686 -115 -682
rect 126 -657 130 -653
rect 138 -664 142 -660
rect 169 -653 173 -649
rect 297 -645 301 -641
rect 309 -652 313 -648
rect 340 -641 344 -637
rect 536 -631 540 -627
rect 570 -635 574 -631
rect 582 -642 586 -638
rect 613 -631 617 -627
rect 51 -700 55 -696
rect 17 -716 21 -712
rect 63 -703 67 -699
rect 94 -696 98 -692
rect 789 -696 793 -692
rect 140 -745 144 -741
rect 297 -734 301 -730
rect 148 -752 152 -748
rect 176 -759 180 -755
rect 309 -741 313 -737
rect 321 -748 325 -744
rect 333 -755 337 -751
rect 358 -730 362 -726
rect -206 -786 -202 -782
rect -194 -793 -190 -789
rect -168 -786 -164 -782
rect -131 -786 -127 -782
rect -156 -801 -152 -797
rect -97 -786 -93 -782
rect -119 -793 -115 -789
rect 17 -776 21 -772
rect 51 -780 55 -776
rect 63 -787 67 -783
rect 94 -776 98 -772
rect 570 -722 574 -718
rect 536 -738 540 -734
rect 582 -725 586 -721
rect 613 -718 617 -714
rect 801 -703 805 -699
rect 827 -696 831 -692
rect 864 -696 868 -692
rect 839 -711 843 -707
rect 898 -696 902 -692
rect 876 -703 880 -699
rect 398 -773 402 -769
rect 129 -819 133 -815
rect 141 -826 145 -822
rect 172 -815 176 -811
rect 406 -780 410 -776
rect 414 -787 418 -783
rect 659 -767 663 -763
rect 457 -780 461 -776
rect 667 -774 671 -770
rect 695 -781 699 -777
rect 422 -794 426 -790
rect 536 -798 540 -794
rect 570 -802 574 -798
rect 582 -809 586 -805
rect 613 -798 617 -794
rect 297 -832 301 -828
rect 51 -862 55 -858
rect -206 -893 -202 -889
rect -194 -900 -190 -896
rect -168 -893 -164 -889
rect -131 -893 -127 -889
rect -156 -908 -152 -904
rect -97 -893 -93 -889
rect -119 -900 -115 -896
rect 17 -878 21 -874
rect 63 -865 67 -861
rect 94 -858 98 -854
rect 309 -839 313 -835
rect 321 -846 325 -842
rect 351 -828 355 -824
rect 789 -803 793 -799
rect 801 -810 805 -806
rect 827 -803 831 -799
rect 864 -803 868 -799
rect 839 -818 843 -814
rect 898 -803 902 -799
rect 876 -810 880 -806
rect 571 -887 575 -883
rect 137 -907 141 -903
rect 537 -903 541 -899
rect 583 -890 587 -886
rect 614 -883 618 -879
rect 145 -914 149 -910
rect 173 -921 177 -917
rect 17 -938 21 -934
rect 51 -942 55 -938
rect 63 -949 67 -945
rect 94 -938 98 -934
rect 297 -925 301 -921
rect 309 -932 313 -928
rect 340 -921 344 -917
rect 789 -910 793 -906
rect 660 -932 664 -928
rect 668 -939 672 -935
rect 696 -946 700 -942
rect 801 -917 805 -913
rect 827 -910 831 -906
rect 864 -910 868 -906
rect 839 -925 843 -921
rect 898 -910 902 -906
rect 876 -917 880 -913
rect 537 -963 541 -959
rect -206 -1000 -202 -996
rect -194 -1007 -190 -1003
rect -168 -1000 -164 -996
rect -131 -1000 -127 -996
rect -156 -1015 -152 -1011
rect -97 -1000 -93 -996
rect -119 -1007 -115 -1003
rect 126 -981 130 -977
rect 138 -988 142 -984
rect 169 -977 173 -973
rect 571 -967 575 -963
rect 583 -974 587 -970
rect 614 -963 618 -959
rect -206 -1107 -202 -1103
rect -194 -1114 -190 -1110
rect -168 -1107 -164 -1103
rect -131 -1107 -127 -1103
rect -156 -1122 -152 -1118
rect -97 -1107 -93 -1103
rect -119 -1114 -115 -1110
<< polypplus >>
rect -164 -240 -162 -228
rect -127 -240 -125 -228
rect -164 -347 -162 -335
rect -127 -347 -125 -335
rect -164 -454 -162 -442
rect -127 -454 -125 -442
rect 831 -471 833 -459
rect 868 -471 870 -459
rect -164 -561 -162 -549
rect -127 -561 -125 -549
rect 831 -578 833 -566
rect 868 -578 870 -566
rect -164 -668 -162 -656
rect -127 -668 -125 -656
rect 831 -685 833 -673
rect -164 -775 -162 -763
rect -127 -775 -125 -763
rect 868 -685 870 -673
rect -164 -882 -162 -870
rect -127 -882 -125 -870
rect 831 -792 833 -780
rect 868 -792 870 -780
rect 831 -899 833 -887
rect 868 -899 870 -887
rect -164 -989 -162 -977
rect -127 -989 -125 -977
rect -164 -1096 -162 -1084
rect -127 -1096 -125 -1084
<< metal1 >>
rect -209 -212 -91 -207
rect -209 -216 -205 -212
rect -171 -216 -167 -212
rect -134 -216 -130 -212
rect -98 -216 -94 -212
rect -210 -251 -206 -247
rect -185 -262 -181 -240
rect -147 -247 -143 -228
rect -110 -247 -106 -228
rect -90 -247 -86 -228
rect -147 -251 -131 -247
rect -110 -251 -97 -247
rect -90 -251 200 -247
rect -185 -266 -156 -262
rect -185 -278 -181 -266
rect -147 -272 -143 -251
rect -110 -272 -106 -251
rect -90 -278 -86 -251
rect -209 -288 -205 -284
rect -171 -288 -167 -284
rect -134 -288 -130 -284
rect -98 -288 -94 -284
rect -209 -293 -91 -288
rect -209 -319 -91 -314
rect -209 -323 -205 -319
rect -171 -323 -167 -319
rect -134 -323 -130 -319
rect -98 -323 -94 -319
rect -210 -358 -206 -354
rect -185 -369 -181 -347
rect -147 -354 -143 -335
rect -110 -354 -106 -335
rect -90 -354 -86 -335
rect 44 -345 94 -341
rect 50 -349 54 -345
rect 70 -349 74 -345
rect -147 -358 -131 -354
rect -110 -358 -97 -354
rect -90 -358 -82 -354
rect -185 -373 -156 -369
rect -185 -385 -181 -373
rect -147 -379 -143 -358
rect -110 -379 -106 -358
rect -90 -385 -86 -358
rect 10 -363 34 -359
rect 90 -349 94 -345
rect 16 -367 20 -363
rect 60 -368 64 -361
rect 60 -372 94 -368
rect 104 -370 108 -361
rect 24 -388 28 -379
rect 38 -376 51 -372
rect 38 -388 42 -376
rect 59 -381 63 -375
rect 52 -385 63 -381
rect 72 -388 76 -372
rect -209 -395 -205 -391
rect -171 -395 -167 -391
rect -134 -395 -130 -391
rect -98 -395 -94 -391
rect -3 -392 17 -388
rect 24 -392 42 -388
rect 24 -395 28 -392
rect -209 -400 -91 -395
rect 104 -374 126 -370
rect 104 -394 108 -374
rect 16 -405 20 -401
rect 47 -405 51 -400
rect 90 -405 94 -400
rect 10 -409 34 -405
rect 44 -409 94 -405
rect 122 -417 126 -374
rect 129 -380 168 -376
rect 135 -384 139 -380
rect 164 -402 168 -380
rect 164 -406 179 -402
rect -209 -426 -91 -421
rect 10 -423 34 -419
rect 44 -423 94 -419
rect 122 -421 140 -417
rect -209 -430 -205 -426
rect -171 -430 -167 -426
rect -134 -430 -130 -426
rect -98 -430 -94 -426
rect 16 -427 20 -423
rect 50 -427 54 -423
rect 70 -427 74 -423
rect 90 -427 94 -423
rect -210 -465 -206 -461
rect -185 -476 -181 -454
rect -147 -461 -143 -442
rect -110 -461 -106 -442
rect -90 -461 -86 -442
rect 24 -448 28 -439
rect 60 -448 64 -439
rect 104 -448 108 -439
rect 122 -428 148 -424
rect 122 -448 126 -428
rect 155 -431 159 -408
rect 175 -410 179 -406
rect 196 -411 200 -251
rect 563 -360 613 -356
rect 569 -364 573 -360
rect 589 -364 593 -360
rect 529 -378 553 -374
rect 609 -364 613 -360
rect 535 -382 539 -378
rect 579 -383 583 -376
rect 579 -387 613 -383
rect 623 -385 627 -376
rect 543 -403 547 -394
rect 557 -391 570 -387
rect 557 -403 561 -391
rect 578 -396 582 -390
rect 571 -400 582 -396
rect 591 -403 595 -387
rect 516 -407 536 -403
rect 543 -407 561 -403
rect 543 -410 547 -407
rect 196 -415 484 -411
rect 623 -389 645 -385
rect 623 -409 627 -389
rect 183 -431 187 -422
rect 283 -423 502 -419
rect 535 -420 539 -416
rect 566 -420 570 -415
rect 609 -420 613 -415
rect 283 -431 287 -423
rect 290 -430 340 -426
rect 370 -430 409 -426
rect 145 -435 176 -431
rect 183 -435 287 -431
rect 296 -434 300 -430
rect 316 -434 320 -430
rect 145 -438 149 -435
rect 183 -438 187 -435
rect 135 -448 139 -444
rect 155 -448 159 -444
rect 175 -448 179 -444
rect 336 -434 340 -430
rect 376 -434 380 -430
rect 6 -452 17 -448
rect 24 -452 46 -448
rect 60 -452 94 -448
rect 104 -452 126 -448
rect 129 -452 179 -448
rect 24 -455 28 -452
rect -147 -465 -131 -461
rect -110 -465 -97 -461
rect -90 -465 -82 -461
rect 42 -456 51 -452
rect 16 -465 20 -461
rect 39 -463 63 -459
rect -185 -480 -156 -476
rect -185 -492 -181 -480
rect -147 -486 -143 -465
rect -110 -486 -106 -465
rect -90 -492 -86 -465
rect 10 -469 34 -465
rect 1 -489 5 -470
rect 39 -480 43 -463
rect 72 -466 76 -452
rect 104 -472 108 -452
rect 306 -455 310 -446
rect 350 -455 354 -446
rect 122 -462 172 -458
rect 306 -459 340 -455
rect 350 -459 367 -455
rect 405 -452 409 -430
rect 405 -456 420 -452
rect 128 -466 132 -462
rect 148 -466 152 -462
rect 168 -466 172 -462
rect 242 -463 297 -459
rect 47 -483 51 -478
rect 90 -483 94 -478
rect 44 -486 94 -483
rect 138 -487 142 -478
rect 182 -487 186 -478
rect 242 -487 246 -463
rect 1 -491 109 -489
rect 138 -491 172 -487
rect 182 -491 246 -487
rect 1 -493 129 -491
rect 105 -495 129 -493
rect -209 -502 -205 -498
rect -171 -502 -167 -498
rect -134 -502 -130 -498
rect -98 -502 -94 -498
rect -3 -498 102 -496
rect -3 -500 141 -498
rect 98 -502 141 -500
rect -209 -507 -91 -502
rect 44 -507 94 -503
rect 150 -505 154 -491
rect 50 -511 54 -507
rect 70 -511 74 -507
rect 10 -525 34 -521
rect 90 -511 94 -507
rect 182 -511 186 -491
rect 125 -522 129 -517
rect 168 -522 172 -517
rect -209 -533 -91 -528
rect 16 -529 20 -525
rect -209 -537 -205 -533
rect -171 -537 -167 -533
rect -134 -537 -130 -533
rect -98 -537 -94 -533
rect 60 -530 64 -523
rect 60 -534 94 -530
rect 104 -532 108 -523
rect 122 -526 172 -522
rect -210 -572 -206 -568
rect -185 -583 -181 -561
rect -147 -568 -143 -549
rect -110 -568 -106 -549
rect -90 -568 -86 -549
rect 24 -550 28 -541
rect 38 -538 51 -534
rect 38 -550 42 -538
rect 59 -543 63 -537
rect 52 -547 63 -543
rect 72 -550 76 -534
rect -3 -554 17 -550
rect 24 -554 42 -550
rect 24 -557 28 -554
rect 104 -536 123 -532
rect 104 -556 108 -536
rect 16 -567 20 -563
rect 47 -567 51 -562
rect 90 -567 94 -562
rect -147 -572 -131 -568
rect -110 -572 -97 -568
rect -90 -572 -82 -568
rect 10 -571 34 -567
rect 44 -571 94 -567
rect -185 -587 -156 -583
rect -185 -599 -181 -587
rect -147 -593 -143 -572
rect -110 -593 -106 -572
rect -90 -599 -86 -572
rect 119 -579 123 -536
rect 126 -542 165 -538
rect 132 -546 136 -542
rect 161 -564 165 -542
rect 242 -560 246 -491
rect 259 -470 309 -466
rect 259 -550 263 -470
rect 318 -473 322 -459
rect 350 -479 354 -459
rect 363 -467 367 -459
rect 363 -471 381 -467
rect 363 -478 389 -474
rect 293 -490 297 -485
rect 336 -490 340 -485
rect 290 -494 340 -490
rect 363 -497 367 -478
rect 396 -481 400 -458
rect 416 -460 420 -456
rect 424 -481 428 -472
rect 498 -472 502 -423
rect 529 -424 553 -420
rect 563 -424 613 -420
rect 641 -432 645 -389
rect 648 -395 687 -391
rect 654 -399 658 -395
rect 683 -417 687 -395
rect 683 -421 698 -417
rect 529 -438 553 -434
rect 563 -438 613 -434
rect 641 -436 659 -432
rect 535 -442 539 -438
rect 569 -442 573 -438
rect 589 -442 593 -438
rect 609 -442 613 -438
rect 543 -463 547 -454
rect 579 -463 583 -454
rect 623 -463 627 -454
rect 641 -443 667 -439
rect 641 -463 645 -443
rect 674 -446 678 -423
rect 694 -425 698 -421
rect 702 -446 706 -437
rect 786 -443 904 -438
rect 664 -450 695 -446
rect 702 -450 767 -446
rect 664 -453 668 -450
rect 702 -453 706 -450
rect 654 -463 658 -459
rect 674 -463 678 -459
rect 694 -463 698 -459
rect 525 -467 536 -463
rect 543 -467 565 -463
rect 579 -467 613 -463
rect 623 -467 645 -463
rect 648 -467 698 -463
rect 529 -472 532 -467
rect 543 -470 547 -467
rect 498 -476 532 -472
rect 561 -471 570 -467
rect 535 -480 539 -476
rect 558 -478 582 -474
rect 386 -485 417 -481
rect 424 -485 500 -481
rect 529 -484 553 -480
rect 386 -488 390 -485
rect 424 -488 428 -485
rect 267 -501 367 -497
rect 376 -498 380 -494
rect 396 -498 400 -494
rect 416 -498 420 -494
rect 267 -541 271 -501
rect 370 -502 420 -498
rect 290 -517 351 -513
rect 296 -521 300 -517
rect 318 -521 322 -517
rect 347 -521 351 -517
rect 306 -542 310 -533
rect 328 -542 332 -533
rect 361 -542 365 -533
rect 306 -546 351 -542
rect 361 -546 384 -542
rect 264 -553 277 -550
rect 264 -554 309 -553
rect 273 -557 309 -554
rect 242 -564 321 -560
rect 161 -568 176 -564
rect 10 -585 34 -581
rect 44 -585 94 -581
rect 119 -583 137 -579
rect 16 -589 20 -585
rect 50 -589 54 -585
rect 70 -589 74 -585
rect 90 -589 94 -585
rect -209 -609 -205 -605
rect -171 -609 -167 -605
rect -134 -609 -130 -605
rect -98 -609 -94 -605
rect -209 -614 -91 -609
rect 24 -610 28 -601
rect 60 -610 64 -601
rect 104 -610 108 -601
rect 119 -590 145 -586
rect 119 -610 123 -590
rect 152 -593 156 -570
rect 172 -572 176 -568
rect 180 -593 184 -584
rect 142 -597 173 -593
rect 180 -597 233 -593
rect 142 -600 146 -597
rect 180 -600 184 -597
rect 132 -610 136 -606
rect 152 -610 156 -606
rect 172 -610 176 -606
rect 6 -614 17 -610
rect 24 -614 46 -610
rect 60 -614 94 -610
rect 104 -614 123 -610
rect 126 -614 176 -610
rect 24 -617 28 -614
rect 42 -618 51 -614
rect 16 -627 20 -623
rect 39 -625 63 -621
rect 10 -631 34 -627
rect -209 -640 -91 -635
rect -209 -644 -205 -640
rect -171 -644 -167 -640
rect -134 -644 -130 -640
rect -98 -644 -94 -640
rect 1 -651 5 -632
rect 39 -642 43 -625
rect 72 -628 76 -614
rect 104 -634 108 -614
rect 119 -624 169 -620
rect 125 -628 129 -624
rect 145 -628 149 -624
rect 165 -628 169 -624
rect 47 -645 51 -640
rect 90 -645 94 -640
rect 44 -648 94 -645
rect 135 -649 139 -640
rect 179 -649 183 -640
rect 1 -653 109 -651
rect 135 -653 169 -649
rect 179 -653 232 -649
rect 1 -655 126 -653
rect -210 -679 -206 -675
rect -185 -690 -181 -668
rect -147 -675 -143 -656
rect -110 -675 -106 -656
rect -90 -675 -86 -656
rect 105 -657 126 -655
rect -3 -660 102 -658
rect -3 -662 138 -660
rect 98 -664 138 -662
rect 44 -669 94 -665
rect 147 -667 151 -653
rect 50 -673 54 -669
rect 70 -673 74 -669
rect -147 -679 -131 -675
rect -110 -679 -97 -675
rect -90 -679 -82 -675
rect -185 -694 -156 -690
rect -185 -706 -181 -694
rect -147 -700 -143 -679
rect -110 -700 -106 -679
rect -90 -706 -86 -679
rect 10 -687 34 -683
rect 90 -673 94 -669
rect 179 -673 183 -653
rect 122 -684 126 -679
rect 165 -684 169 -679
rect 16 -691 20 -687
rect 60 -692 64 -685
rect 60 -696 94 -692
rect 104 -694 108 -685
rect 119 -688 169 -684
rect 24 -712 28 -703
rect 38 -700 51 -696
rect 38 -712 42 -700
rect 59 -705 63 -699
rect 52 -709 63 -705
rect 72 -712 76 -696
rect -209 -716 -205 -712
rect -171 -716 -167 -712
rect -134 -716 -130 -712
rect -98 -716 -94 -712
rect -209 -721 -91 -716
rect -3 -716 17 -712
rect 24 -716 42 -712
rect 24 -719 28 -716
rect 104 -698 126 -694
rect 104 -718 108 -698
rect 16 -729 20 -725
rect 47 -729 51 -724
rect 90 -729 94 -724
rect 10 -733 34 -729
rect 44 -733 94 -729
rect 122 -741 126 -698
rect 129 -704 168 -700
rect 135 -708 139 -704
rect 164 -726 168 -704
rect 164 -730 179 -726
rect -209 -747 -91 -742
rect 10 -747 34 -743
rect 44 -747 94 -743
rect 122 -745 140 -741
rect -209 -751 -205 -747
rect -171 -751 -167 -747
rect -134 -751 -130 -747
rect -98 -751 -94 -747
rect 16 -751 20 -747
rect 50 -751 54 -747
rect 70 -751 74 -747
rect 90 -751 94 -747
rect -210 -786 -206 -782
rect -185 -797 -181 -775
rect -147 -782 -143 -763
rect -110 -782 -106 -763
rect -90 -782 -86 -763
rect 24 -772 28 -763
rect 60 -772 64 -763
rect 104 -772 108 -763
rect 122 -752 148 -748
rect 122 -772 126 -752
rect 155 -755 159 -732
rect 175 -734 179 -730
rect 242 -751 246 -564
rect 328 -567 332 -546
rect 259 -593 263 -574
rect 255 -597 263 -593
rect 259 -744 263 -597
rect 268 -648 272 -573
rect 361 -570 365 -546
rect 293 -584 297 -579
rect 347 -584 351 -576
rect 290 -588 351 -584
rect 380 -585 384 -546
rect 387 -548 432 -544
rect 393 -552 397 -548
rect 428 -556 432 -548
rect 428 -560 446 -556
rect 442 -564 446 -560
rect 421 -585 425 -576
rect 450 -585 454 -576
rect 380 -589 398 -585
rect 421 -589 443 -585
rect 450 -589 493 -585
rect 363 -596 406 -592
rect 290 -612 340 -608
rect 296 -616 300 -612
rect 316 -616 320 -612
rect 336 -616 340 -612
rect 306 -637 310 -628
rect 350 -637 354 -628
rect 363 -637 367 -596
rect 276 -648 280 -640
rect 306 -641 340 -637
rect 350 -641 367 -637
rect 379 -603 414 -599
rect 268 -652 309 -648
rect 268 -731 272 -652
rect 318 -655 322 -641
rect 350 -661 354 -641
rect 293 -672 297 -667
rect 336 -672 340 -667
rect 290 -676 340 -672
rect 379 -679 383 -603
rect 421 -606 425 -589
rect 450 -592 454 -589
rect 442 -602 446 -598
rect 403 -610 425 -606
rect 403 -613 407 -610
rect 421 -613 425 -610
rect 428 -606 446 -602
rect 393 -623 397 -619
rect 411 -623 415 -619
rect 428 -623 432 -606
rect 387 -627 432 -623
rect 276 -683 383 -679
rect 276 -714 280 -683
rect 290 -701 358 -697
rect 296 -705 300 -701
rect 318 -705 322 -701
rect 340 -705 344 -701
rect 354 -705 358 -701
rect 306 -726 310 -717
rect 330 -726 334 -717
rect 368 -726 372 -717
rect 306 -730 358 -726
rect 368 -730 384 -726
rect 277 -734 297 -730
rect 259 -748 321 -744
rect 242 -755 333 -751
rect 145 -759 176 -755
rect 340 -758 344 -730
rect 145 -762 149 -759
rect 135 -772 139 -768
rect 155 -772 159 -768
rect 175 -772 179 -768
rect 6 -776 17 -772
rect 24 -776 46 -772
rect 60 -776 94 -772
rect 104 -776 126 -772
rect 129 -776 179 -772
rect 24 -779 28 -776
rect -147 -786 -131 -782
rect -110 -786 -97 -782
rect -90 -786 -82 -782
rect 42 -780 51 -776
rect -185 -801 -156 -797
rect -185 -813 -181 -801
rect -147 -807 -143 -786
rect -110 -807 -106 -786
rect -90 -813 -86 -786
rect 16 -789 20 -785
rect 39 -787 63 -783
rect 10 -793 34 -789
rect 1 -813 5 -794
rect 39 -804 43 -787
rect 72 -790 76 -776
rect 104 -796 108 -776
rect 122 -786 172 -782
rect 128 -790 132 -786
rect 148 -790 152 -786
rect 168 -790 172 -786
rect 47 -807 51 -802
rect 90 -807 94 -802
rect 44 -810 94 -807
rect 138 -811 142 -802
rect 182 -811 186 -802
rect 255 -811 259 -764
rect 1 -815 109 -813
rect 138 -815 172 -811
rect 182 -815 259 -811
rect 1 -817 129 -815
rect 105 -819 129 -817
rect -209 -823 -205 -819
rect -171 -823 -167 -819
rect -134 -823 -130 -819
rect -98 -823 -94 -819
rect -209 -828 -91 -823
rect -3 -822 102 -820
rect -3 -824 141 -822
rect 98 -826 141 -824
rect 44 -831 94 -827
rect 150 -829 154 -815
rect 50 -835 54 -831
rect 70 -835 74 -831
rect 10 -849 34 -845
rect 90 -835 94 -831
rect 182 -835 186 -815
rect 125 -846 129 -841
rect 168 -846 172 -841
rect -209 -854 -91 -849
rect 16 -853 20 -849
rect -209 -858 -205 -854
rect -171 -858 -167 -854
rect -134 -858 -130 -854
rect -98 -858 -94 -854
rect 60 -854 64 -847
rect 60 -858 94 -854
rect 104 -856 108 -847
rect 122 -850 172 -846
rect -210 -893 -206 -889
rect -185 -904 -181 -882
rect -147 -889 -143 -870
rect -110 -889 -106 -870
rect -90 -889 -86 -870
rect 24 -874 28 -865
rect 38 -862 51 -858
rect 38 -874 42 -862
rect 59 -867 63 -861
rect 52 -871 63 -867
rect 72 -874 76 -858
rect -3 -878 17 -874
rect 24 -878 42 -874
rect 24 -881 28 -878
rect 104 -860 123 -856
rect 104 -880 108 -860
rect -147 -893 -131 -889
rect -110 -893 -97 -889
rect -90 -893 -82 -889
rect 16 -891 20 -887
rect 47 -891 51 -886
rect 90 -891 94 -886
rect -185 -908 -156 -904
rect -185 -920 -181 -908
rect -147 -914 -143 -893
rect -110 -914 -106 -893
rect -90 -920 -86 -893
rect 10 -895 34 -891
rect 44 -895 94 -891
rect 119 -903 123 -860
rect 126 -866 165 -862
rect 132 -870 136 -866
rect 161 -888 165 -866
rect 161 -892 176 -888
rect 10 -909 34 -905
rect 44 -909 94 -905
rect 119 -907 137 -903
rect 16 -913 20 -909
rect 50 -913 54 -909
rect 70 -913 74 -909
rect 90 -913 94 -909
rect -209 -930 -205 -926
rect -171 -930 -167 -926
rect -134 -930 -130 -926
rect -98 -930 -94 -926
rect -209 -935 -91 -930
rect 24 -934 28 -925
rect 60 -934 64 -925
rect 104 -934 108 -925
rect 119 -914 145 -910
rect 119 -934 123 -914
rect 152 -917 156 -894
rect 172 -896 176 -892
rect 180 -917 184 -908
rect 142 -921 173 -917
rect 180 -921 246 -917
rect 142 -924 146 -921
rect 180 -924 184 -921
rect 132 -934 136 -930
rect 152 -934 156 -930
rect 255 -928 259 -815
rect 267 -842 271 -764
rect 276 -828 280 -764
rect 368 -761 372 -730
rect 293 -775 297 -770
rect 354 -775 358 -767
rect 380 -769 384 -730
rect 387 -732 441 -728
rect 393 -736 397 -732
rect 437 -747 441 -732
rect 437 -751 460 -747
rect 380 -773 398 -769
rect 290 -779 358 -775
rect 429 -776 433 -760
rect 456 -755 460 -751
rect 464 -776 468 -767
rect 475 -776 479 -680
rect 373 -780 406 -776
rect 429 -780 457 -776
rect 464 -780 479 -776
rect 290 -799 351 -795
rect 296 -803 300 -799
rect 318 -803 322 -799
rect 347 -803 351 -799
rect 306 -824 310 -815
rect 328 -824 332 -815
rect 361 -824 365 -815
rect 373 -824 377 -780
rect 306 -828 351 -824
rect 361 -828 377 -824
rect 380 -794 422 -790
rect 276 -832 297 -828
rect 276 -833 280 -832
rect 267 -846 321 -842
rect 328 -849 332 -828
rect 275 -917 279 -855
rect 361 -852 365 -828
rect 293 -866 297 -861
rect 347 -866 351 -858
rect 290 -870 351 -866
rect 290 -892 340 -888
rect 296 -896 300 -892
rect 316 -896 320 -892
rect 336 -896 340 -892
rect 268 -921 279 -917
rect 306 -917 310 -908
rect 350 -917 354 -908
rect 380 -917 384 -794
rect 429 -798 433 -780
rect 464 -783 468 -780
rect 456 -793 460 -789
rect 403 -802 433 -798
rect 442 -797 460 -793
rect 403 -805 407 -802
rect 419 -805 423 -802
rect 393 -815 397 -811
rect 411 -815 415 -811
rect 429 -815 433 -811
rect 442 -815 446 -797
rect 387 -819 446 -815
rect 489 -891 493 -589
rect 496 -726 500 -485
rect 558 -495 562 -478
rect 591 -481 595 -467
rect 623 -487 627 -467
rect 763 -478 767 -450
rect 786 -447 790 -443
rect 824 -447 828 -443
rect 861 -447 865 -443
rect 897 -447 901 -443
rect 763 -482 789 -478
rect 810 -493 814 -471
rect 848 -478 852 -459
rect 885 -478 889 -459
rect 905 -478 909 -459
rect 848 -482 864 -478
rect 885 -482 898 -478
rect 905 -482 913 -478
rect 566 -498 570 -493
rect 609 -498 613 -493
rect 563 -502 613 -498
rect 810 -497 839 -493
rect 810 -509 814 -497
rect 848 -503 852 -482
rect 885 -503 889 -482
rect 905 -509 909 -482
rect 786 -519 790 -515
rect 824 -519 828 -515
rect 861 -519 865 -515
rect 897 -519 901 -515
rect 563 -524 613 -520
rect 786 -524 904 -519
rect 569 -528 573 -524
rect 589 -528 593 -524
rect 529 -542 553 -538
rect 609 -528 613 -524
rect 535 -546 539 -542
rect 579 -547 583 -540
rect 579 -551 613 -547
rect 623 -549 627 -540
rect 543 -567 547 -558
rect 557 -555 570 -551
rect 557 -567 561 -555
rect 578 -560 582 -554
rect 571 -564 582 -560
rect 591 -567 595 -551
rect 516 -571 536 -567
rect 543 -571 561 -567
rect 543 -574 547 -571
rect 623 -553 645 -549
rect 623 -573 627 -553
rect 535 -584 539 -580
rect 566 -584 570 -579
rect 609 -584 613 -579
rect 529 -588 553 -584
rect 563 -588 613 -584
rect 641 -596 645 -553
rect 786 -550 904 -545
rect 786 -554 790 -550
rect 824 -554 828 -550
rect 861 -554 865 -550
rect 897 -554 901 -550
rect 648 -559 687 -555
rect 654 -563 658 -559
rect 683 -581 687 -559
rect 683 -585 698 -581
rect 529 -602 553 -598
rect 563 -602 613 -598
rect 641 -600 659 -596
rect 535 -606 539 -602
rect 569 -606 573 -602
rect 589 -606 593 -602
rect 609 -606 613 -602
rect 543 -627 547 -618
rect 579 -627 583 -618
rect 623 -627 627 -618
rect 641 -607 667 -603
rect 641 -627 645 -607
rect 674 -610 678 -587
rect 694 -589 698 -585
rect 763 -589 789 -585
rect 702 -610 706 -601
rect 763 -610 767 -589
rect 664 -614 695 -610
rect 702 -614 767 -610
rect 810 -600 814 -578
rect 848 -585 852 -566
rect 885 -585 889 -566
rect 905 -585 909 -566
rect 848 -589 864 -585
rect 885 -589 898 -585
rect 905 -589 913 -585
rect 810 -604 839 -600
rect 664 -617 668 -614
rect 702 -617 706 -614
rect 810 -616 814 -604
rect 848 -610 852 -589
rect 885 -610 889 -589
rect 654 -627 658 -623
rect 674 -627 678 -623
rect 905 -616 909 -589
rect 694 -627 698 -623
rect 525 -631 536 -627
rect 543 -631 565 -627
rect 579 -631 613 -627
rect 623 -631 645 -627
rect 648 -631 698 -627
rect 786 -626 790 -622
rect 824 -626 828 -622
rect 861 -626 865 -622
rect 897 -626 901 -622
rect 786 -631 904 -626
rect 543 -634 547 -631
rect 561 -635 570 -631
rect 535 -644 539 -640
rect 558 -642 582 -638
rect 529 -648 553 -644
rect 558 -659 562 -642
rect 591 -645 595 -631
rect 623 -651 627 -631
rect 786 -657 904 -652
rect 566 -662 570 -657
rect 609 -662 613 -657
rect 563 -665 613 -662
rect 786 -661 790 -657
rect 824 -661 828 -657
rect 861 -661 865 -657
rect 897 -661 901 -657
rect 509 -679 767 -675
rect 563 -691 613 -687
rect 569 -695 573 -691
rect 589 -695 593 -691
rect 529 -709 553 -705
rect 609 -695 613 -691
rect 763 -692 767 -679
rect 763 -696 789 -692
rect 535 -713 539 -709
rect 579 -714 583 -707
rect 579 -718 613 -714
rect 623 -716 627 -707
rect 810 -707 814 -685
rect 848 -692 852 -673
rect 885 -692 889 -673
rect 905 -692 909 -673
rect 848 -696 864 -692
rect 885 -696 898 -692
rect 905 -696 913 -692
rect 810 -711 839 -707
rect 496 -730 529 -726
rect 525 -734 529 -730
rect 543 -734 547 -725
rect 557 -722 570 -718
rect 557 -734 561 -722
rect 578 -727 582 -721
rect 571 -731 582 -727
rect 591 -734 595 -718
rect 516 -738 536 -734
rect 543 -738 561 -734
rect 543 -741 547 -738
rect 623 -720 645 -716
rect 623 -740 627 -720
rect 535 -751 539 -747
rect 566 -751 570 -746
rect 609 -751 613 -746
rect 529 -755 553 -751
rect 563 -755 613 -751
rect 641 -763 645 -720
rect 648 -726 687 -722
rect 810 -723 814 -711
rect 848 -717 852 -696
rect 885 -717 889 -696
rect 654 -730 658 -726
rect 683 -748 687 -726
rect 905 -723 909 -696
rect 786 -733 790 -729
rect 824 -733 828 -729
rect 861 -733 865 -729
rect 897 -733 901 -729
rect 786 -738 904 -733
rect 683 -752 698 -748
rect 529 -769 553 -765
rect 563 -769 613 -765
rect 641 -767 659 -763
rect 535 -773 539 -769
rect 569 -773 573 -769
rect 589 -773 593 -769
rect 609 -773 613 -769
rect 543 -794 547 -785
rect 579 -794 583 -785
rect 623 -794 627 -785
rect 641 -774 667 -770
rect 641 -794 645 -774
rect 674 -777 678 -754
rect 694 -756 698 -752
rect 702 -777 706 -768
rect 786 -764 904 -759
rect 786 -768 790 -764
rect 824 -768 828 -764
rect 861 -768 865 -764
rect 897 -768 901 -764
rect 664 -781 695 -777
rect 702 -781 767 -777
rect 664 -784 668 -781
rect 702 -784 706 -781
rect 654 -794 658 -790
rect 674 -794 678 -790
rect 694 -794 698 -790
rect 525 -798 536 -794
rect 543 -798 565 -794
rect 579 -798 613 -794
rect 623 -798 645 -794
rect 648 -798 698 -794
rect 543 -801 547 -798
rect 561 -802 570 -798
rect 535 -811 539 -807
rect 558 -809 582 -805
rect 529 -815 553 -811
rect 558 -826 562 -809
rect 591 -812 595 -798
rect 623 -818 627 -798
rect 763 -799 767 -781
rect 763 -803 789 -799
rect 810 -814 814 -792
rect 848 -799 852 -780
rect 885 -799 889 -780
rect 905 -799 909 -780
rect 848 -803 864 -799
rect 885 -803 898 -799
rect 905 -803 913 -799
rect 810 -818 839 -814
rect 566 -829 570 -824
rect 609 -829 613 -824
rect 563 -832 613 -829
rect 810 -830 814 -818
rect 848 -824 852 -803
rect 885 -824 889 -803
rect 905 -830 909 -803
rect 786 -840 790 -836
rect 824 -840 828 -836
rect 861 -840 865 -836
rect 897 -840 901 -836
rect 786 -845 904 -840
rect 564 -856 614 -852
rect 570 -860 574 -856
rect 590 -860 594 -856
rect 530 -874 554 -870
rect 610 -860 614 -856
rect 536 -878 540 -874
rect 580 -879 584 -872
rect 580 -883 614 -879
rect 624 -881 628 -872
rect 786 -871 904 -866
rect 786 -875 790 -871
rect 824 -875 828 -871
rect 861 -875 865 -871
rect 897 -875 901 -871
rect 489 -895 530 -891
rect 526 -899 530 -895
rect 544 -899 548 -890
rect 558 -887 571 -883
rect 558 -899 562 -887
rect 579 -892 583 -886
rect 572 -896 583 -892
rect 592 -899 596 -883
rect 517 -903 537 -899
rect 544 -903 562 -899
rect 544 -906 548 -903
rect 624 -885 646 -881
rect 624 -905 628 -885
rect 536 -916 540 -912
rect 567 -916 571 -911
rect 610 -916 614 -911
rect 306 -921 340 -917
rect 350 -921 384 -917
rect 530 -920 554 -916
rect 564 -920 614 -916
rect 275 -925 297 -921
rect 172 -934 176 -930
rect 255 -932 309 -928
rect 6 -938 17 -934
rect 24 -938 46 -934
rect 60 -938 94 -934
rect 104 -938 123 -934
rect 126 -938 176 -934
rect 318 -935 322 -921
rect 24 -941 28 -938
rect 42 -942 51 -938
rect 16 -951 20 -947
rect 39 -949 63 -945
rect 10 -955 34 -951
rect -209 -961 -91 -956
rect -209 -965 -205 -961
rect -171 -965 -167 -961
rect -134 -965 -130 -961
rect -98 -965 -94 -961
rect -210 -1000 -206 -996
rect -185 -1011 -181 -989
rect -147 -996 -143 -977
rect -110 -996 -106 -977
rect -90 -996 -86 -977
rect 1 -975 5 -956
rect 39 -966 43 -949
rect 72 -952 76 -938
rect 104 -958 108 -938
rect 119 -948 169 -944
rect 125 -952 129 -948
rect 145 -952 149 -948
rect 165 -952 169 -948
rect 350 -941 354 -921
rect 642 -928 646 -885
rect 649 -891 688 -887
rect 655 -895 659 -891
rect 684 -913 688 -891
rect 763 -910 789 -906
rect 684 -917 699 -913
rect 530 -934 554 -930
rect 564 -934 614 -930
rect 642 -932 660 -928
rect 536 -938 540 -934
rect 570 -938 574 -934
rect 590 -938 594 -934
rect 293 -952 297 -947
rect 336 -952 340 -947
rect 610 -938 614 -934
rect 290 -956 340 -952
rect 544 -959 548 -950
rect 580 -959 584 -950
rect 624 -959 628 -950
rect 642 -939 668 -935
rect 642 -959 646 -939
rect 675 -942 679 -919
rect 695 -921 699 -917
rect 703 -942 707 -933
rect 763 -942 767 -910
rect 810 -921 814 -899
rect 848 -906 852 -887
rect 885 -906 889 -887
rect 905 -906 909 -887
rect 848 -910 864 -906
rect 885 -910 898 -906
rect 905 -910 913 -906
rect 810 -925 839 -921
rect 810 -937 814 -925
rect 848 -931 852 -910
rect 885 -931 889 -910
rect 665 -946 696 -942
rect 703 -946 767 -942
rect 905 -937 909 -910
rect 665 -949 669 -946
rect 703 -949 707 -946
rect 655 -959 659 -955
rect 675 -959 679 -955
rect 786 -947 790 -943
rect 824 -947 828 -943
rect 861 -947 865 -943
rect 897 -947 901 -943
rect 786 -952 904 -947
rect 695 -959 699 -955
rect 526 -963 537 -959
rect 544 -963 566 -959
rect 580 -963 614 -959
rect 624 -963 646 -959
rect 649 -963 699 -959
rect 47 -969 51 -964
rect 90 -969 94 -964
rect 44 -972 94 -969
rect 135 -973 139 -964
rect 544 -966 548 -963
rect 562 -967 571 -963
rect 1 -977 109 -975
rect 135 -977 169 -973
rect 536 -976 540 -972
rect 559 -974 583 -970
rect 1 -979 126 -977
rect 105 -981 126 -979
rect -3 -984 102 -982
rect -3 -986 138 -984
rect 98 -988 138 -986
rect 147 -991 151 -977
rect 530 -980 554 -976
rect 559 -991 563 -974
rect 592 -977 596 -963
rect 624 -983 628 -963
rect -147 -1000 -131 -996
rect -110 -1000 -97 -996
rect -90 -1000 -82 -996
rect -185 -1015 -156 -1011
rect -185 -1027 -181 -1015
rect -147 -1021 -143 -1000
rect -110 -1021 -106 -1000
rect -90 -1027 -86 -1000
rect 567 -994 571 -989
rect 610 -994 614 -989
rect 564 -998 614 -994
rect 122 -1008 126 -1003
rect 165 -1008 169 -1003
rect 119 -1012 169 -1008
rect -209 -1037 -205 -1033
rect -171 -1037 -167 -1033
rect -134 -1037 -130 -1033
rect -98 -1037 -94 -1033
rect -209 -1042 -91 -1037
rect -209 -1068 -91 -1063
rect -209 -1072 -205 -1068
rect -171 -1072 -167 -1068
rect -134 -1072 -130 -1068
rect -98 -1072 -94 -1068
rect -210 -1107 -206 -1103
rect -185 -1118 -181 -1096
rect -147 -1103 -143 -1084
rect -110 -1103 -106 -1084
rect -90 -1103 -86 -1084
rect -147 -1107 -131 -1103
rect -110 -1107 -97 -1103
rect -90 -1107 -82 -1103
rect -185 -1122 -156 -1118
rect -185 -1134 -181 -1122
rect -147 -1128 -143 -1107
rect -110 -1128 -106 -1107
rect -90 -1134 -86 -1107
rect -209 -1144 -205 -1140
rect -171 -1144 -167 -1140
rect -134 -1144 -130 -1140
rect -98 -1144 -94 -1140
rect -209 -1149 -91 -1144
<< m2contact >>
rect -82 -358 -77 -353
rect 47 -385 52 -380
rect -8 -393 -3 -388
rect 566 -400 571 -395
rect 511 -408 516 -403
rect 484 -415 489 -410
rect 1 -453 6 -448
rect -82 -465 -77 -460
rect 1 -470 6 -465
rect 34 -480 39 -475
rect -8 -500 -3 -495
rect 47 -547 52 -542
rect -8 -555 -3 -550
rect -82 -572 -77 -567
rect 254 -498 259 -493
rect 246 -515 251 -510
rect 520 -468 525 -463
rect 267 -546 272 -541
rect 259 -555 264 -550
rect 233 -597 238 -592
rect 1 -615 6 -610
rect 1 -632 6 -627
rect 34 -642 39 -637
rect 232 -653 237 -648
rect -8 -662 -3 -657
rect -82 -679 -77 -674
rect 47 -709 52 -704
rect -8 -717 -3 -712
rect 259 -574 264 -569
rect 268 -573 273 -568
rect 250 -597 255 -592
rect 276 -640 281 -635
rect 475 -680 480 -675
rect 276 -719 281 -714
rect 267 -736 272 -731
rect 276 -739 281 -734
rect 255 -764 260 -759
rect 266 -764 271 -759
rect 1 -777 6 -772
rect -82 -786 -77 -781
rect 1 -794 6 -789
rect 34 -804 39 -799
rect -8 -824 -3 -819
rect 47 -871 52 -866
rect -8 -879 -3 -874
rect -82 -893 -77 -888
rect 246 -921 251 -916
rect 276 -764 281 -759
rect 275 -838 280 -833
rect 275 -855 280 -850
rect 263 -921 268 -916
rect 279 -880 284 -875
rect 553 -495 558 -490
rect 566 -564 571 -559
rect 511 -572 516 -567
rect 520 -632 525 -627
rect 553 -659 558 -654
rect 504 -680 509 -675
rect 566 -731 571 -726
rect 511 -739 516 -734
rect 520 -799 525 -794
rect 553 -826 558 -821
rect 567 -896 572 -891
rect 512 -904 517 -899
rect 1 -939 6 -934
rect 1 -956 6 -951
rect 34 -966 39 -961
rect 521 -964 526 -959
rect -8 -986 -3 -981
rect 554 -991 559 -986
rect -82 -1000 -77 -995
rect -82 -1107 -77 -1102
<< metal2 >>
rect -198 -251 -168 -247
rect -198 -254 -194 -251
rect -221 -258 -194 -254
rect -172 -254 -168 -251
rect -172 -258 -119 -254
rect -221 -301 -217 -258
rect -221 -305 759 -301
rect -221 -361 -217 -305
rect -198 -358 -168 -354
rect 1 -354 41 -352
rect -77 -356 41 -354
rect -77 -358 5 -356
rect -198 -361 -194 -358
rect -221 -365 -194 -361
rect -172 -361 -168 -358
rect -172 -365 -119 -361
rect -221 -468 -217 -365
rect -198 -465 -168 -461
rect -8 -461 -4 -393
rect -77 -465 -4 -461
rect -198 -468 -194 -465
rect -221 -472 -194 -468
rect -172 -468 -168 -465
rect -172 -472 -119 -468
rect -221 -575 -217 -472
rect -8 -476 -4 -465
rect 1 -448 5 -358
rect 37 -368 41 -356
rect 37 -371 47 -368
rect 43 -385 47 -371
rect 520 -371 560 -367
rect 511 -411 515 -408
rect 489 -415 515 -411
rect 1 -465 5 -453
rect -8 -480 34 -476
rect -8 -495 -4 -480
rect 511 -491 515 -415
rect 520 -463 524 -371
rect 556 -383 560 -371
rect 556 -386 566 -383
rect 562 -400 566 -386
rect 755 -485 759 -305
rect 797 -482 827 -478
rect 797 -485 801 -482
rect 755 -489 801 -485
rect 823 -485 827 -482
rect 823 -489 876 -485
rect 511 -495 553 -491
rect 254 -502 257 -498
rect 254 -506 543 -502
rect 1 -518 41 -514
rect 251 -514 507 -510
rect 1 -542 5 -518
rect 37 -530 41 -518
rect 37 -533 47 -530
rect -17 -546 5 -542
rect -198 -572 -168 -568
rect -17 -568 -13 -546
rect -77 -572 -13 -568
rect -198 -575 -194 -572
rect -221 -579 -194 -575
rect -172 -575 -168 -572
rect -172 -579 -119 -575
rect -221 -682 -217 -579
rect -8 -638 -4 -555
rect 1 -610 5 -546
rect 43 -547 47 -533
rect 259 -569 263 -555
rect 268 -568 272 -546
rect 288 -550 297 -546
rect 238 -597 250 -593
rect 1 -627 5 -615
rect -8 -642 34 -638
rect 255 -640 276 -636
rect -8 -651 -4 -642
rect -16 -655 -4 -651
rect 255 -649 259 -640
rect 237 -653 259 -649
rect 288 -641 292 -550
rect 503 -576 507 -514
rect 539 -531 543 -506
rect 520 -535 560 -531
rect 511 -576 515 -572
rect 503 -580 515 -576
rect 288 -645 297 -641
rect -198 -679 -168 -675
rect -16 -675 -12 -655
rect -8 -657 -4 -655
rect -77 -679 -12 -675
rect -198 -682 -194 -679
rect -221 -686 -194 -682
rect -172 -682 -168 -679
rect 1 -680 41 -676
rect -172 -686 -119 -682
rect -221 -789 -217 -686
rect 1 -704 5 -680
rect 37 -692 41 -680
rect 288 -692 292 -645
rect 511 -655 515 -580
rect 520 -627 524 -535
rect 556 -547 560 -535
rect 556 -550 566 -547
rect 562 -564 566 -550
rect 755 -592 759 -489
rect 797 -589 827 -585
rect 797 -592 801 -589
rect 755 -596 801 -592
rect 823 -592 827 -589
rect 823 -596 876 -592
rect 511 -659 553 -655
rect 480 -679 504 -675
rect 37 -695 47 -692
rect -16 -708 5 -704
rect -198 -786 -168 -782
rect -16 -782 -12 -708
rect -77 -786 -12 -782
rect -198 -789 -194 -786
rect -221 -793 -194 -789
rect -172 -789 -168 -786
rect -172 -793 -119 -789
rect -221 -896 -217 -793
rect -8 -800 -4 -717
rect 1 -772 5 -708
rect 43 -709 47 -695
rect 288 -696 524 -692
rect 276 -723 280 -719
rect 255 -727 280 -723
rect 183 -755 187 -746
rect 183 -759 251 -755
rect 183 -762 187 -759
rect 247 -768 251 -759
rect 255 -759 259 -727
rect 267 -759 271 -736
rect 277 -759 281 -739
rect 288 -737 292 -696
rect 520 -698 524 -696
rect 520 -702 560 -698
rect 288 -741 309 -737
rect 288 -768 292 -741
rect 247 -772 292 -768
rect 1 -789 5 -777
rect 190 -787 246 -783
rect -8 -804 34 -800
rect -8 -811 -4 -804
rect -16 -815 -4 -811
rect -16 -858 -12 -815
rect -8 -819 -4 -815
rect -73 -862 -12 -858
rect 1 -842 41 -838
rect -198 -893 -168 -889
rect -73 -889 -69 -862
rect 1 -866 5 -842
rect 37 -854 41 -842
rect 37 -857 47 -854
rect -77 -893 -69 -889
rect -16 -870 5 -866
rect -198 -896 -194 -893
rect -221 -900 -194 -896
rect -172 -896 -168 -893
rect -172 -900 -119 -896
rect -221 -1003 -217 -900
rect -16 -954 -12 -870
rect -73 -958 -12 -954
rect -198 -1000 -168 -996
rect -73 -996 -69 -958
rect -8 -962 -4 -879
rect 1 -934 5 -870
rect 43 -871 47 -857
rect 1 -951 5 -939
rect -8 -966 34 -962
rect -8 -973 -4 -966
rect -77 -1000 -69 -996
rect -16 -977 -4 -973
rect -198 -1003 -194 -1000
rect -221 -1007 -194 -1003
rect -172 -1003 -168 -1000
rect -172 -1007 -119 -1003
rect -221 -1110 -217 -1007
rect -198 -1107 -168 -1103
rect -16 -1103 -12 -977
rect -8 -981 -4 -977
rect 179 -973 183 -964
rect 190 -973 194 -787
rect 288 -835 292 -772
rect 305 -787 414 -783
rect 511 -822 515 -739
rect 520 -794 524 -702
rect 556 -714 560 -702
rect 755 -699 759 -596
rect 797 -696 827 -692
rect 797 -699 801 -696
rect 755 -703 801 -699
rect 823 -699 827 -696
rect 823 -703 876 -699
rect 556 -717 566 -714
rect 562 -731 566 -717
rect 755 -806 759 -703
rect 797 -803 827 -799
rect 797 -806 801 -803
rect 755 -810 801 -806
rect 823 -806 827 -803
rect 823 -810 876 -806
rect 511 -826 553 -822
rect 275 -850 279 -838
rect 288 -839 309 -835
rect 521 -867 561 -863
rect 521 -875 525 -867
rect 284 -879 525 -875
rect 251 -921 263 -917
rect 179 -977 194 -973
rect 179 -997 183 -977
rect 512 -987 516 -904
rect 521 -959 525 -879
rect 557 -879 561 -867
rect 557 -882 567 -879
rect 563 -896 567 -882
rect 755 -913 759 -810
rect 797 -910 827 -906
rect 797 -913 801 -910
rect 755 -917 801 -913
rect 823 -913 827 -910
rect 823 -917 876 -913
rect 512 -991 554 -987
rect -77 -1107 -12 -1103
rect -198 -1110 -194 -1107
rect -221 -1114 -194 -1110
rect -172 -1110 -168 -1107
rect -172 -1114 -119 -1110
<< m3contact >>
rect 246 -788 251 -783
rect 300 -788 305 -783
<< metal3 >>
rect 251 -787 300 -783
<< labels >>
rlabel metal1 537 -377 537 -377 5 VDD
rlabel metal1 540 -422 540 -422 1 GND
rlabel metal1 537 -437 537 -437 5 VDD
rlabel metal1 540 -482 540 -482 1 GND
rlabel metal1 581 -436 581 -436 5 VDD
rlabel metal1 595 -500 595 -500 1 GND
rlabel metal1 581 -358 581 -358 5 VDD
rlabel metal1 595 -422 595 -422 1 GND
rlabel metal1 665 -393 665 -393 5 VDD
rlabel metal1 666 -465 666 -465 1 GND
rlabel ndcontact 537 -413 537 -413 1 GND
rlabel pdcontact 537 -388 537 -388 1 VDD
rlabel ndcontact 568 -409 568 -409 1 GND
rlabel pdcontact 571 -370 571 -370 1 VDD
rlabel pdcontact 591 -370 591 -370 1 VDD
rlabel pdcontact 611 -370 611 -370 1 VDD
rlabel ndcontact 611 -412 611 -412 1 GND
rlabel ndcontact 656 -456 656 -456 1 GND
rlabel ndcontact 676 -456 676 -456 1 GND
rlabel ndcontact 696 -456 696 -456 1 GND
rlabel pdcontact 696 -431 696 -431 1 VDD
rlabel pdcontact 696 -762 696 -762 1 VDD
rlabel ndcontact 696 -787 696 -787 1 GND
rlabel ndcontact 676 -787 676 -787 1 GND
rlabel ndcontact 656 -787 656 -787 1 GND
rlabel ndcontact 611 -821 611 -821 1 GND
rlabel pdcontact 611 -779 611 -779 1 VDD
rlabel ndcontact 611 -743 611 -743 1 GND
rlabel pdcontact 611 -701 611 -701 1 VDD
rlabel pdcontact 591 -701 591 -701 1 VDD
rlabel pdcontact 571 -701 571 -701 1 VDD
rlabel ndcontact 568 -740 568 -740 1 GND
rlabel pdcontact 591 -779 591 -779 1 VDD
rlabel pdcontact 571 -779 571 -779 1 VDD
rlabel ndcontact 568 -818 568 -818 1 GND
rlabel pdcontact 537 -719 537 -719 1 VDD
rlabel ndcontact 537 -744 537 -744 1 GND
rlabel pdcontact 537 -779 537 -779 1 VDD
rlabel ndcontact 537 -804 537 -804 1 GND
rlabel metal1 666 -796 666 -796 1 GND
rlabel metal1 665 -724 665 -724 5 VDD
rlabel metal1 595 -753 595 -753 1 GND
rlabel metal1 581 -689 581 -689 5 VDD
rlabel metal1 595 -831 595 -831 1 GND
rlabel metal1 581 -767 581 -767 5 VDD
rlabel metal1 540 -813 540 -813 1 GND
rlabel metal1 537 -768 537 -768 5 VDD
rlabel metal1 540 -753 540 -753 1 GND
rlabel metal1 537 -708 537 -708 5 VDD
rlabel metal1 537 -541 537 -541 5 VDD
rlabel metal1 540 -586 540 -586 1 GND
rlabel metal1 537 -601 537 -601 5 VDD
rlabel metal1 540 -646 540 -646 1 GND
rlabel metal1 581 -600 581 -600 5 VDD
rlabel metal1 595 -664 595 -664 1 GND
rlabel metal1 581 -522 581 -522 5 VDD
rlabel metal1 595 -586 595 -586 1 GND
rlabel metal1 665 -557 665 -557 5 VDD
rlabel metal1 666 -629 666 -629 1 GND
rlabel ndcontact 537 -637 537 -637 1 GND
rlabel pdcontact 537 -612 537 -612 1 VDD
rlabel ndcontact 537 -577 537 -577 1 GND
rlabel pdcontact 537 -552 537 -552 1 VDD
rlabel ndcontact 568 -651 568 -651 1 GND
rlabel pdcontact 571 -612 571 -612 1 VDD
rlabel pdcontact 591 -612 591 -612 1 VDD
rlabel ndcontact 568 -573 568 -573 1 GND
rlabel pdcontact 571 -534 571 -534 1 VDD
rlabel pdcontact 591 -534 591 -534 1 VDD
rlabel pdcontact 611 -534 611 -534 1 VDD
rlabel ndcontact 611 -576 611 -576 1 GND
rlabel pdcontact 611 -612 611 -612 1 VDD
rlabel ndcontact 611 -654 611 -654 1 GND
rlabel ndcontact 656 -620 656 -620 1 GND
rlabel ndcontact 676 -620 676 -620 1 GND
rlabel ndcontact 696 -620 696 -620 1 GND
rlabel pdcontact 696 -595 696 -595 1 VDD
rlabel metal1 538 -873 538 -873 5 VDD
rlabel metal1 541 -918 541 -918 1 GND
rlabel metal1 538 -933 538 -933 5 VDD
rlabel metal1 541 -978 541 -978 1 GND
rlabel metal1 582 -932 582 -932 5 VDD
rlabel metal1 596 -996 596 -996 1 GND
rlabel metal1 582 -854 582 -854 5 VDD
rlabel metal1 596 -918 596 -918 1 GND
rlabel metal1 666 -889 666 -889 5 VDD
rlabel metal1 667 -961 667 -961 1 GND
rlabel ndcontact 538 -969 538 -969 1 GND
rlabel pdcontact 538 -944 538 -944 1 VDD
rlabel ndcontact 538 -909 538 -909 1 GND
rlabel pdcontact 538 -884 538 -884 1 VDD
rlabel ndcontact 569 -983 569 -983 1 GND
rlabel pdcontact 572 -944 572 -944 1 VDD
rlabel pdcontact 592 -944 592 -944 1 VDD
rlabel ndcontact 569 -905 569 -905 1 GND
rlabel pdcontact 572 -866 572 -866 1 VDD
rlabel pdcontact 592 -866 592 -866 1 VDD
rlabel pdcontact 612 -866 612 -866 1 VDD
rlabel ndcontact 612 -908 612 -908 1 GND
rlabel pdcontact 612 -944 612 -944 1 VDD
rlabel ndcontact 612 -986 612 -986 1 GND
rlabel ndcontact 657 -952 657 -952 1 GND
rlabel ndcontact 677 -952 677 -952 1 GND
rlabel ndcontact 697 -952 697 -952 1 GND
rlabel pdcontact 697 -927 697 -927 1 VDD
rlabel polycontact 538 -465 538 -465 1 p0
rlabel pdcontact 545 -448 545 -448 1 p0_bar
rlabel polycontact 572 -469 572 -469 1 p0_bar
rlabel polycontact 584 -476 584 -476 1 c0
rlabel polycontact 538 -405 538 -405 1 c0
rlabel pdcontact 545 -388 545 -388 1 c0_bar
rlabel polycontact 572 -389 572 -389 1 c0_bar
rlabel polycontact 584 -392 584 -392 1 p0
rlabel metal1 708 -448 708 -448 7 s0
rlabel ndcontact 704 -456 704 -456 1 s0
rlabel pdcontact 704 -431 704 -431 1 s0
rlabel pdcontact 656 -411 656 -411 1 vdd
rlabel pdcontact 581 -370 581 -370 1 a1n
rlabel ndiffusion 581 -409 581 -409 1 a1m
rlabel ndcontact 593 -409 593 -409 1 a1n
rlabel polycontact 615 -385 615 -385 1 a1n
rlabel ndcontact 625 -412 625 -412 1 outa1
rlabel pdcontact 625 -370 625 -370 1 outa1
rlabel polycontact 661 -434 661 -434 1 outa1
rlabel polycontact 669 -441 669 -441 1 outa2
rlabel polycontact 697 -448 697 -448 1 s0_bar
rlabel ndcontact 666 -456 666 -456 1 s0_bar
rlabel pdcontact 676 -411 676 -411 1 s0_bar
rlabel pdcontact 625 -448 625 -448 1 outa2
rlabel ndcontact 625 -490 625 -490 1 outa2
rlabel polycontact 615 -465 615 -465 1 a2n
rlabel pdcontact 581 -448 581 -448 1 a2n
rlabel ndcontact 593 -487 593 -487 1 a2n
rlabel ndiffusion 581 -487 581 -487 1 a2m
rlabel polycontact 538 -629 538 -629 1 p1
rlabel ndcontact 545 -637 545 -637 1 p1_bar
rlabel pdcontact 545 -612 545 -612 1 p1_bar
rlabel polycontact 572 -633 572 -633 1 p1_bar
rlabel pdcontact 581 -612 581 -612 1 b2n
rlabel ndcontact 593 -651 593 -651 1 b2n
rlabel ndiffusion 581 -651 581 -651 1 b2m
rlabel polycontact 615 -629 615 -629 1 b2n
rlabel pdcontact 625 -612 625 -612 1 outb2
rlabel ndcontact 625 -654 625 -654 1 outb2
rlabel polycontact 669 -605 669 -605 1 outb2
rlabel ndcontact 666 -620 666 -620 1 s1_bar
rlabel polycontact 697 -612 697 -612 1 s1_bar
rlabel metal1 708 -612 708 -612 7 s1
rlabel ndcontact 704 -620 704 -620 1 s1
rlabel pdcontact 704 -595 704 -595 1 s1
rlabel pdcontact 676 -575 676 -575 1 s1_bar
rlabel pdcontact 656 -575 656 -575 1 vdd
rlabel polycontact 661 -598 661 -598 1 outb1
rlabel ndcontact 625 -576 625 -576 1 outb1
rlabel pdcontact 625 -534 625 -534 1 outb1
rlabel polycontact 615 -549 615 -549 1 b1n
rlabel pdcontact 581 -534 581 -534 1 b1n
rlabel ndcontact 593 -573 593 -573 1 b1n
rlabel ndiffusion 581 -573 581 -573 1 b1m
rlabel polycontact 584 -556 584 -556 1 p1
rlabel polycontact 572 -553 572 -553 1 c1_bar
rlabel ndcontact 545 -577 545 -577 1 c1_bar
rlabel pdcontact 545 -552 545 -552 1 c1_bar
rlabel polycontact 538 -796 538 -796 1 p2
rlabel ndcontact 545 -804 545 -804 1 p2_bar
rlabel pdcontact 545 -779 545 -779 1 p2_bar
rlabel polycontact 572 -800 572 -800 1 p2_bar
rlabel polycontact 584 -807 584 -807 1 c2
rlabel polycontact 538 -736 538 -736 1 c2
rlabel polycontact 584 -723 584 -723 1 p2
rlabel pdcontact 581 -701 581 -701 1 c1n
rlabel ndcontact 593 -740 593 -740 1 c1n
rlabel ndiffusion 581 -740 581 -740 1 c1m
rlabel polycontact 615 -716 615 -716 1 c1n
rlabel pdcontact 625 -701 625 -701 1 outc1
rlabel ndcontact 625 -743 625 -743 1 outc1
rlabel polycontact 661 -765 661 -765 1 outc1
rlabel pdcontact 656 -742 656 -742 1 vdd
rlabel polycontact 669 -772 669 -772 1 outc2
rlabel pdcontact 676 -742 676 -742 1 s2_bar
rlabel polycontact 697 -779 697 -779 1 s2_bar
rlabel ndcontact 666 -787 666 -787 1 s2_bar
rlabel metal1 708 -779 708 -779 7 s2
rlabel pdcontact 581 -779 581 -779 1 c2n
rlabel ndiffusion 581 -818 581 -818 1 c2m
rlabel ndcontact 593 -818 593 -818 1 c2n
rlabel polycontact 615 -796 615 -796 1 c2n
rlabel ndcontact 625 -821 625 -821 1 outc2
rlabel pdcontact 625 -779 625 -779 1 outc2
rlabel polycontact 539 -961 539 -961 1 p3
rlabel ndcontact 546 -969 546 -969 1 p3_bar
rlabel pdcontact 546 -944 546 -944 1 p3_bar
rlabel polycontact 573 -965 573 -965 1 p3_bar
rlabel polycontact 585 -972 585 -972 1 c3
rlabel polycontact 539 -901 539 -901 1 c3
rlabel polycontact 585 -888 585 -888 1 p3
rlabel pdcontact 582 -866 582 -866 1 d1n
rlabel ndcontact 594 -905 594 -905 1 d1n
rlabel ndiffusion 582 -905 582 -905 1 d1m
rlabel polycontact 616 -881 616 -881 1 d1n
rlabel pdcontact 626 -866 626 -866 1 outd1
rlabel ndcontact 626 -908 626 -908 1 outd1
rlabel polycontact 662 -930 662 -930 1 outd1
rlabel polycontact 670 -937 670 -937 1 outd2
rlabel pdcontact 657 -907 657 -907 1 vdd
rlabel pdcontact 677 -907 677 -907 1 s3_bar
rlabel polycontact 698 -944 698 -944 1 s3_bar
rlabel metal1 709 -944 709 -944 7 s3
rlabel pdcontact 705 -927 705 -927 1 s3
rlabel ndcontact 667 -952 667 -952 1 s3_bar
rlabel pdcontact 582 -944 582 -944 1 d2n
rlabel ndcontact 594 -983 594 -983 1 d2n
rlabel ndiffusion 582 -983 582 -983 1 d2m
rlabel polycontact 616 -961 616 -961 1 d2n
rlabel pdcontact 626 -944 626 -944 1 outd2
rlabel ndcontact 626 -986 626 -986 1 outd2
rlabel pdiffusion 667 -906 667 -906 1 dps
rlabel pdiffusion 666 -742 666 -742 1 cps
rlabel pdiffusion 666 -574 666 -574 1 bps
rlabel pdiffusion 666 -412 666 -412 1 aps
rlabel ndcontact 704 -787 704 -787 1 s2
rlabel pdcontact 704 -762 704 -762 1 s2
rlabel ndcontact 705 -952 705 -952 1 s3
rlabel ndcontact 545 -413 545 -413 1 c0_bar
rlabel ndcontact 545 -473 545 -473 1 p0_bar
rlabel pdcontact 537 -448 537 -448 1 vdd
rlabel ndcontact 537 -473 537 -473 1 gnd
rlabel ndcontact 568 -487 568 -487 1 gnd
rlabel pdcontact 571 -448 571 -448 1 vdd
rlabel pdcontact 591 -448 591 -448 1 vdd
rlabel ndcontact 611 -490 611 -490 1 gnd
rlabel pdcontact 611 -448 611 -448 1 vdd
rlabel metal1 404 -730 404 -730 5 VDD
rlabel pdcontact 395 -748 395 -748 1 vdd
rlabel metal1 405 -817 405 -817 1 GND
rlabel ndcontact 413 -808 413 -808 1 gnd
rlabel ndcontact 395 -808 395 -808 1 gnd
rlabel ndcontact 431 -808 431 -808 1 gnd
rlabel ndcontact 458 -786 458 -786 1 gnd
rlabel pdcontact 458 -761 458 -761 1 vdd
rlabel metal1 308 -797 308 -797 5 VDD
rlabel metal1 295 -868 295 -868 2 GND
rlabel ndcontact 295 -855 295 -855 3 gnd
rlabel ndcontact 349 -855 349 -855 1 gnd
rlabel pdcontact 349 -809 349 -809 1 vdd
rlabel pdcontact 320 -809 320 -809 1 vdd
rlabel pdcontact 298 -809 298 -809 1 vdd
rlabel metal1 308 -428 308 -428 5 VDD
rlabel metal1 295 -492 295 -492 2 GND
rlabel metal1 388 -500 388 -500 1 GND
rlabel metal1 387 -428 387 -428 5 VDD
rlabel metal1 308 -515 308 -515 5 VDD
rlabel metal1 295 -586 295 -586 2 GND
rlabel ndcontact 295 -573 295 -573 3 gnd
rlabel ndcontact 349 -573 349 -573 1 gnd
rlabel pdcontact 349 -527 349 -527 1 vdd
rlabel pdcontact 320 -527 320 -527 1 vdd
rlabel pdcontact 298 -527 298 -527 1 vdd
rlabel metal1 308 -610 308 -610 5 VDD
rlabel metal1 295 -674 295 -674 2 GND
rlabel metal1 404 -546 404 -546 5 VDD
rlabel metal1 405 -625 405 -625 1 GND
rlabel ndcontact 444 -595 444 -595 1 gnd
rlabel pdcontact 444 -570 444 -570 1 vdd
rlabel ndcontact 413 -616 413 -616 1 gnd
rlabel ndcontact 395 -616 395 -616 1 gnd
rlabel pdcontact 395 -564 395 -564 1 vdd
rlabel metal1 308 -699 308 -699 5 VDD
rlabel pdcontact 320 -711 320 -711 1 vdd
rlabel pdcontact 298 -711 298 -711 1 vdd
rlabel ndcontact 295 -764 295 -764 3 gnd
rlabel metal1 295 -777 295 -777 2 GND
rlabel pdcontact 356 -711 356 -711 1 vdd
rlabel ndcontact 356 -764 356 -764 1 gnd
rlabel pdcontact 342 -711 342 -711 1 vdd
rlabel metal1 308 -890 308 -890 5 VDD
rlabel metal1 295 -954 295 -954 2 GND
rlabel polycontact 299 -461 299 -461 1 g0
rlabel polycontact 342 -457 342 -457 1 p1g0_bar
rlabel polycontact 383 -469 383 -469 1 p1g0
rlabel polycontact 391 -476 391 -476 1 g1
rlabel polycontact 419 -483 419 -483 1 c2_bar
rlabel metal1 430 -483 430 -483 1 c2
rlabel pdcontact 298 -440 298 -440 1 vdd
rlabel pdcontact 318 -440 318 -440 1 vdd
rlabel pdcontact 308 -440 308 -440 1 p1g0_bar
rlabel ndcontact 320 -479 320 -479 1 p1g0_bar
rlabel ndcontact 295 -479 295 -479 3 gnd
rlabel pdcontact 338 -440 338 -440 1 vdd
rlabel pdcontact 352 -440 352 -440 1 p1g0
rlabel ndcontact 338 -482 338 -482 1 gnd
rlabel ndcontact 352 -482 352 -482 1 p1g0
rlabel pdcontact 378 -446 378 -446 1 vdd
rlabel ndcontact 378 -491 378 -491 1 gnd
rlabel ndcontact 398 -491 398 -491 1 gnd
rlabel ndcontact 388 -491 388 -491 1 c2_bar
rlabel pdcontact 398 -446 398 -446 1 c2_bar
rlabel ndcontact 418 -491 418 -491 1 gnd
rlabel ndcontact 426 -491 426 -491 1 c2
rlabel pdcontact 426 -466 426 -466 1 c2
rlabel pdcontact 418 -466 418 -466 1 vdd
rlabel ndiffusion 308 -479 308 -479 1 n1
rlabel pdiffusion 388 -445 388 -445 1 n2
rlabel polycontact 323 -562 323 -562 1 g0
rlabel ndiffusion 308 -573 308 -573 1 n3
rlabel ndiffusion 320 -573 320 -573 1 n4
rlabel polycontact 353 -544 353 -544 1 p2p1g0_bar
rlabel pdcontact 330 -527 330 -527 1 p2p1g0_bar
rlabel pdcontact 308 -527 308 -527 1 p2p1g0_bar
rlabel pdcontact 363 -527 363 -527 1 p2p1g0
rlabel ndcontact 363 -573 363 -573 1 p2p1g0
rlabel ndcontact 330 -573 330 -573 1 p2p1g0_bar
rlabel polycontact 400 -587 400 -587 1 p2p1g0
rlabel pdcontact 318 -622 318 -622 1 vdd
rlabel pdcontact 338 -622 338 -622 1 vdd
rlabel pdcontact 298 -622 298 -622 1 vdd
rlabel polycontact 311 -650 311 -650 1 g1
rlabel polycontact 342 -639 342 -639 1 p2g1_bar
rlabel pdcontact 308 -622 308 -622 1 p2g1_bar
rlabel ndcontact 320 -661 320 -661 1 p2g1_bar
rlabel ndcontact 295 -661 295 -661 3 gnd
rlabel ndcontact 338 -664 338 -664 1 gnd
rlabel pdcontact 352 -622 352 -622 1 p2g1
rlabel ndcontact 352 -664 352 -664 1 p2g1
rlabel polycontact 408 -594 408 -594 1 p2g1
rlabel polycontact 416 -601 416 -601 1 g2
rlabel ndcontact 452 -595 452 -595 1 c3
rlabel pdcontact 452 -570 452 -570 1 c3
rlabel polycontact 335 -753 335 -753 1 g0
rlabel ndiffusion 308 -661 308 -661 1 n5
rlabel pdiffusion 405 -564 405 -564 1 n6
rlabel pdiffusion 413 -564 413 -564 1 n7
rlabel ndiffusion 308 -764 308 -764 1 n8
rlabel ndiffusion 320 -764 320 -764 1 n9
rlabel ndiffusion 332 -764 332 -764 1 n10
rlabel ndcontact 342 -764 342 -764 1 p3p2p1g0_bar
rlabel pdcontact 332 -711 332 -711 1 p3p2p1g0_bar
rlabel pdcontact 308 -711 308 -711 1 p3p2p1g0_bar
rlabel polycontact 360 -728 360 -728 1 p3p2p1g0_bar
rlabel ndcontact 370 -764 370 -764 1 p3p2p1g0
rlabel pdcontact 370 -711 370 -711 1 p3p2p1g0
rlabel polycontact 400 -771 400 -771 1 p3p2p1g0
rlabel polycontact 323 -844 323 -844 1 g1
rlabel ndiffusion 308 -855 308 -855 1 n11
rlabel ndiffusion 320 -855 320 -855 1 n12
rlabel ndcontact 330 -855 330 -855 1 p3p2g1_bar
rlabel pdcontact 308 -809 308 -809 1 p3p2g1_bar
rlabel pdcontact 330 -809 330 -809 1 p3p2g1_bar
rlabel polycontact 353 -826 353 -826 1 p3p2g1_bar
rlabel ndcontact 363 -855 363 -855 1 p3p2g1
rlabel pdcontact 363 -809 363 -809 1 p3p2g1
rlabel polycontact 408 -778 408 -778 1 p3p2g1
rlabel polycontact 311 -930 311 -930 1 g2
rlabel ndcontact 295 -941 295 -941 3 gnd
rlabel ndcontact 338 -944 338 -944 1 gnd
rlabel ndcontact 320 -941 320 -941 1 p3g2_bar
rlabel pdcontact 298 -902 298 -902 1 vdd
rlabel pdcontact 308 -902 308 -902 1 p3g2_bar
rlabel pdcontact 318 -902 318 -902 1 vdd
rlabel polycontact 342 -919 342 -919 1 p3g2_bar
rlabel pdcontact 338 -902 338 -902 1 vdd
rlabel pdcontact 352 -902 352 -902 1 p3g2
rlabel ndcontact 352 -944 352 -944 1 p3g2
rlabel ndiffusion 308 -941 308 -941 1 n13
rlabel polycontact 424 -792 424 -792 1 p3g2
rlabel pdiffusion 405 -747 405 -747 1 n14
rlabel pdiffusion 413 -747 413 -747 1 n15
rlabel pdiffusion 421 -747 421 -747 1 n16
rlabel ndcontact 405 -808 405 -808 1 cout_bar
rlabel ndcontact 421 -808 421 -808 1 cout_bar
rlabel pdcontact 431 -748 431 -748 1 cout_bar
rlabel polycontact 459 -778 459 -778 1 cout_bar
rlabel metal1 470 -778 470 -778 7 cout
rlabel ndcontact 466 -786 466 -786 1 cout
rlabel pdcontact 466 -761 466 -761 1 cout
rlabel polycontact 311 -468 311 -468 1 p1
rlabel polycontact 311 -555 311 -555 1 p1
rlabel polycontact 323 -746 323 -746 1 p1
rlabel polycontact 299 -548 299 -548 1 p2
rlabel polycontact 299 -643 299 -643 1 p2
rlabel polycontact 311 -739 311 -739 1 p2
rlabel polycontact 311 -837 311 -837 1 p2
rlabel polycontact 299 -732 299 -732 1 p3
rlabel polycontact 299 -830 299 -830 1 p3
rlabel polycontact 299 -923 299 -923 1 p3
rlabel metal1 18 -362 18 -362 5 VDD
rlabel metal1 21 -407 21 -407 1 GND
rlabel metal1 18 -422 18 -422 5 VDD
rlabel metal1 21 -467 21 -467 1 GND
rlabel metal1 62 -421 62 -421 5 VDD
rlabel metal1 76 -485 76 -485 1 GND
rlabel metal1 62 -343 62 -343 5 VDD
rlabel metal1 76 -407 76 -407 1 GND
rlabel metal1 146 -378 146 -378 5 VDD
rlabel metal1 147 -450 147 -450 1 GND
rlabel ndcontact 18 -458 18 -458 1 GND
rlabel pdcontact 18 -433 18 -433 1 VDD
rlabel ndcontact 18 -398 18 -398 1 GND
rlabel pdcontact 18 -373 18 -373 1 VDD
rlabel ndcontact 49 -472 49 -472 1 GND
rlabel ndiffusion 62 -472 62 -472 1 and2m
rlabel ndcontact 74 -472 74 -472 1 and2n
rlabel pdcontact 52 -433 52 -433 1 VDD
rlabel pdcontact 62 -433 62 -433 1 and2n
rlabel pdcontact 72 -433 72 -433 1 VDD
rlabel ndcontact 49 -394 49 -394 1 GND
rlabel ndiffusion 62 -394 62 -394 1 and1m
rlabel ndcontact 74 -394 74 -394 1 and1n
rlabel pdcontact 52 -355 52 -355 1 VDD
rlabel pdcontact 72 -355 72 -355 1 VDD
rlabel pdcontact 62 -355 62 -355 1 and1n
rlabel polycontact 96 -370 96 -370 1 and1n
rlabel pdcontact 92 -355 92 -355 1 VDD
rlabel pdcontact 106 -355 106 -355 1 outand1
rlabel ndcontact 106 -397 106 -397 1 outand1
rlabel ndcontact 92 -397 92 -397 1 GND
rlabel pdcontact 92 -433 92 -433 1 VDD
rlabel pdcontact 106 -433 106 -433 1 outand2
rlabel ndcontact 106 -475 106 -475 1 outand2
rlabel ndcontact 92 -475 92 -475 1 GND
rlabel polycontact 96 -450 96 -450 1 and2n
rlabel polycontact 142 -419 142 -419 1 outand1
rlabel polycontact 150 -426 150 -426 1 outand2
rlabel ndcontact 137 -441 137 -441 1 GND
rlabel ndcontact 157 -441 157 -441 1 GND
rlabel ndcontact 177 -441 177 -441 1 GND
rlabel pdcontact 177 -416 177 -416 1 VDD
rlabel metal1 127 -524 127 -524 2 GND
rlabel metal1 140 -460 140 -460 5 VDD
rlabel metal1 18 -524 18 -524 5 VDD
rlabel metal1 21 -569 21 -569 1 GND
rlabel metal1 18 -584 18 -584 5 VDD
rlabel metal1 21 -629 21 -629 1 GND
rlabel metal1 62 -583 62 -583 5 VDD
rlabel metal1 76 -647 76 -647 1 GND
rlabel metal1 62 -505 62 -505 5 VDD
rlabel metal1 76 -569 76 -569 1 GND
rlabel ndcontact 18 -620 18 -620 1 GND
rlabel pdcontact 18 -595 18 -595 1 VDD
rlabel ndcontact 18 -560 18 -560 1 GND
rlabel pdcontact 18 -535 18 -535 1 VDD
rlabel ndcontact 49 -634 49 -634 1 GND
rlabel pdcontact 52 -595 52 -595 1 VDD
rlabel pdcontact 72 -595 72 -595 1 VDD
rlabel ndcontact 49 -556 49 -556 1 GND
rlabel pdcontact 52 -517 52 -517 1 VDD
rlabel pdcontact 72 -517 72 -517 1 VDD
rlabel pdcontact 92 -517 92 -517 1 VDD
rlabel ndcontact 92 -559 92 -559 1 GND
rlabel pdcontact 92 -595 92 -595 1 VDD
rlabel ndcontact 92 -637 92 -637 1 GND
rlabel metal1 143 -540 143 -540 5 VDD
rlabel metal1 144 -612 144 -612 1 GND
rlabel ndcontact 134 -603 134 -603 1 GND
rlabel ndcontact 154 -603 154 -603 1 GND
rlabel ndcontact 174 -603 174 -603 1 GND
rlabel pdcontact 174 -578 174 -578 1 VDD
rlabel metal1 137 -622 137 -622 5 VDD
rlabel metal1 124 -686 124 -686 2 GND
rlabel metal1 18 -686 18 -686 5 VDD
rlabel metal1 21 -731 21 -731 1 GND
rlabel metal1 18 -746 18 -746 5 VDD
rlabel metal1 21 -791 21 -791 1 GND
rlabel metal1 62 -745 62 -745 5 VDD
rlabel metal1 76 -809 76 -809 1 GND
rlabel metal1 62 -667 62 -667 5 VDD
rlabel metal1 76 -731 76 -731 1 GND
rlabel metal1 146 -702 146 -702 5 VDD
rlabel metal1 147 -774 147 -774 1 GND
rlabel ndcontact 18 -782 18 -782 1 GND
rlabel pdcontact 18 -757 18 -757 1 VDD
rlabel ndcontact 18 -722 18 -722 1 GND
rlabel pdcontact 18 -697 18 -697 1 VDD
rlabel ndcontact 49 -796 49 -796 1 GND
rlabel pdcontact 52 -757 52 -757 1 VDD
rlabel pdcontact 72 -757 72 -757 1 VDD
rlabel ndcontact 49 -718 49 -718 1 GND
rlabel pdcontact 52 -679 52 -679 1 VDD
rlabel pdcontact 72 -679 72 -679 1 VDD
rlabel pdcontact 92 -679 92 -679 1 VDD
rlabel ndcontact 92 -721 92 -721 1 GND
rlabel pdcontact 92 -757 92 -757 1 VDD
rlabel ndcontact 92 -799 92 -799 1 GND
rlabel ndcontact 137 -765 137 -765 1 GND
rlabel ndcontact 157 -765 157 -765 1 GND
rlabel ndcontact 177 -765 177 -765 1 GND
rlabel pdcontact 177 -740 177 -740 1 VDD
rlabel metal1 127 -848 127 -848 2 GND
rlabel metal1 140 -784 140 -784 5 VDD
rlabel metal1 18 -848 18 -848 5 VDD
rlabel metal1 21 -893 21 -893 1 GND
rlabel metal1 18 -908 18 -908 5 VDD
rlabel metal1 21 -953 21 -953 1 GND
rlabel metal1 62 -907 62 -907 5 VDD
rlabel metal1 76 -971 76 -971 1 GND
rlabel metal1 62 -829 62 -829 5 VDD
rlabel metal1 76 -893 76 -893 1 GND
rlabel ndcontact 18 -944 18 -944 1 GND
rlabel pdcontact 18 -919 18 -919 1 VDD
rlabel ndcontact 18 -884 18 -884 1 GND
rlabel pdcontact 18 -859 18 -859 1 VDD
rlabel ndcontact 49 -958 49 -958 1 GND
rlabel pdcontact 52 -919 52 -919 1 VDD
rlabel pdcontact 72 -919 72 -919 1 VDD
rlabel ndcontact 49 -880 49 -880 1 GND
rlabel pdcontact 52 -841 52 -841 1 VDD
rlabel pdcontact 72 -841 72 -841 1 VDD
rlabel pdcontact 92 -841 92 -841 1 VDD
rlabel ndcontact 92 -883 92 -883 1 GND
rlabel pdcontact 92 -919 92 -919 1 VDD
rlabel ndcontact 92 -961 92 -961 1 GND
rlabel metal1 143 -864 143 -864 5 VDD
rlabel metal1 144 -936 144 -936 1 GND
rlabel ndcontact 134 -927 134 -927 1 GND
rlabel ndcontact 154 -927 154 -927 1 GND
rlabel ndcontact 174 -927 174 -927 1 GND
rlabel pdcontact 174 -902 174 -902 1 VDD
rlabel metal1 137 -946 137 -946 5 VDD
rlabel metal1 124 -1010 124 -1010 2 GND
rlabel ndcontact 184 -514 184 -514 1 g0
rlabel pdcontact 184 -472 184 -472 1 g0
rlabel ndcontact 170 -514 170 -514 1 gnd
rlabel ndcontact 152 -511 152 -511 1 g0_bar
rlabel polycontact 174 -489 174 -489 1 g0_bar
rlabel pdcontact 140 -472 140 -472 1 g0_bar
rlabel pdcontact 170 -472 170 -472 1 vdd
rlabel pdcontact 150 -472 150 -472 1 vdd
rlabel pdcontact 130 -472 130 -472 1 vdd
rlabel ndcontact 127 -511 127 -511 1 gnd
rlabel ndiffusion 139 -511 139 -511 1 and0m
rlabel polycontact 143 -500 143 -500 1 b0
rlabel ndcontact 185 -441 185 -441 1 p0
rlabel metal1 189 -433 189 -433 7 p0
rlabel pdcontact 185 -416 185 -416 1 p0
rlabel polycontact 178 -433 178 -433 1 p0_bar
rlabel ndcontact 147 -441 147 -441 1 p0_bar
rlabel pdcontact 157 -396 157 -396 1 p0_bar
rlabel pdcontact 137 -396 137 -396 1 vdd
rlabel polycontact 19 -450 19 -450 1 a0
rlabel ndcontact 26 -458 26 -458 1 a0_bar
rlabel pdcontact 26 -433 26 -433 1 a0_bar
rlabel polycontact 53 -454 53 -454 1 a0_bar
rlabel polycontact 65 -461 65 -461 1 b0
rlabel polycontact 19 -390 19 -390 1 b0
rlabel pdcontact 26 -373 26 -373 1 b0_bar
rlabel ndcontact 26 -398 26 -398 1 b0_bar
rlabel polycontact 53 -374 53 -374 1 b0_bar
rlabel polycontact 65 -377 65 -377 1 a0
rlabel polycontact 131 -493 131 -493 1 a0
rlabel ndcontact 167 -676 167 -676 1 gnd
rlabel ndcontact 181 -676 181 -676 1 g1
rlabel pdcontact 181 -634 181 -634 1 g1
rlabel pdcontact 167 -634 167 -634 1 vdd
rlabel polycontact 171 -651 171 -651 1 g1_bar
rlabel ndcontact 149 -673 149 -673 1 g1_bar
rlabel ndcontact 124 -673 124 -673 1 gnd
rlabel pdcontact 137 -634 137 -634 1 g1_bar
rlabel pdcontact 147 -634 147 -634 1 vdd
rlabel pdcontact 127 -634 127 -634 1 vdd
rlabel polycontact 140 -662 140 -662 1 b1
rlabel polycontact 128 -655 128 -655 1 a1
rlabel ndcontact 182 -603 182 -603 1 p1
rlabel pdcontact 182 -578 182 -578 1 p1
rlabel polycontact 175 -595 175 -595 1 p1_bar
rlabel ndcontact 144 -603 144 -603 1 p1_bar
rlabel pdcontact 154 -558 154 -558 1 p1_bar
rlabel pdcontact 134 -558 134 -558 1 vdd
rlabel polycontact 19 -612 19 -612 1 a1
rlabel ndcontact 26 -620 26 -620 1 a1_bar
rlabel pdcontact 26 -595 26 -595 1 a1_bar
rlabel polycontact 53 -616 53 -616 1 a1_bar
rlabel polycontact 65 -623 65 -623 1 b1
rlabel polycontact 19 -552 19 -552 1 b1
rlabel ndcontact 26 -560 26 -560 1 b1_bar
rlabel pdcontact 26 -535 26 -535 1 b1_bar
rlabel polycontact 53 -536 53 -536 1 b1_bar
rlabel polycontact 65 -539 65 -539 1 a1
rlabel metal1 188 -813 188 -813 7 g2
rlabel ndcontact 184 -838 184 -838 1 g2
rlabel pdcontact 184 -796 184 -796 1 g2
rlabel ndcontact 170 -838 170 -838 1 gnd
rlabel ndcontact 152 -835 152 -835 1 g2_bar
rlabel ndcontact 127 -835 127 -835 1 gnd
rlabel polycontact 174 -813 174 -813 1 g2_bar
rlabel polycontact 143 -824 143 -824 1 b2
rlabel polycontact 131 -817 131 -817 1 a2
rlabel pdcontact 170 -796 170 -796 1 vdd
rlabel pdcontact 150 -796 150 -796 1 vdd
rlabel pdcontact 130 -796 130 -796 1 vdd
rlabel pdcontact 140 -796 140 -796 1 g2_bar
rlabel polycontact 178 -757 178 -757 1 p2_bar
rlabel ndcontact 147 -765 147 -765 1 p2_bar
rlabel pdcontact 157 -721 157 -721 1 p2_bar
rlabel pdcontact 137 -720 137 -720 1 vdd
rlabel polycontact 19 -774 19 -774 1 a2
rlabel ndcontact 26 -782 26 -782 1 a2_bar
rlabel pdcontact 26 -757 26 -757 1 a2_bar
rlabel polycontact 53 -778 53 -778 1 a2_bar
rlabel polycontact 65 -785 65 -785 1 b2
rlabel polycontact 19 -714 19 -714 1 b2
rlabel pdcontact 26 -697 26 -697 1 b2_bar
rlabel ndcontact 26 -722 26 -722 1 b2_bar
rlabel polycontact 53 -698 53 -698 1 b2_bar
rlabel polycontact 65 -701 65 -701 1 a2
rlabel ndcontact 167 -1000 167 -1000 1 gnd
rlabel ndcontact 181 -1000 181 -1000 1 g3
rlabel pdcontact 181 -958 181 -958 1 g3
rlabel pdcontact 167 -958 167 -958 1 vdd
rlabel polycontact 171 -975 171 -975 1 g3_bar
rlabel ndcontact 149 -997 149 -997 1 g3_bar
rlabel ndcontact 124 -997 124 -997 1 gnd
rlabel polycontact 140 -986 140 -986 1 b3
rlabel polycontact 128 -979 128 -979 1 a3
rlabel pdcontact 147 -958 147 -958 1 vdd
rlabel pdcontact 127 -958 127 -958 1 vdd
rlabel pdcontact 137 -958 137 -958 1 g3_bar
rlabel ndcontact 182 -927 182 -927 1 p3
rlabel metal1 186 -919 186 -919 1 p3
rlabel pdcontact 182 -902 182 -902 1 p3
rlabel polycontact 175 -919 175 -919 1 p3_bar
rlabel ndcontact 144 -927 144 -927 1 p3_bar
rlabel pdcontact 154 -882 154 -882 1 p3_bar
rlabel pdcontact 134 -882 134 -882 1 vdd
rlabel polycontact 19 -936 19 -936 1 a3
rlabel ndcontact 26 -944 26 -944 1 a3_bar
rlabel pdcontact 26 -919 26 -919 1 a3_bar
rlabel polycontact 53 -940 53 -940 1 a3_bar
rlabel polycontact 65 -947 65 -947 1 b3
rlabel polycontact 19 -876 19 -876 1 b3
rlabel pdcontact 26 -859 26 -859 1 b3_bar
rlabel ndcontact 26 -884 26 -884 1 b3_bar
rlabel polycontact 53 -860 53 -860 1 b3_bar
rlabel polycontact 65 -863 65 -863 1 a3
rlabel polycontact 416 -785 416 -785 1 g3
rlabel pdcontact 185 -740 185 -740 1 p2
rlabel ndcontact 185 -765 185 -765 1 p2
rlabel ndiffusion 62 -556 62 -556 1 anda1m
rlabel ndcontact 74 -556 74 -556 1 anda1n
rlabel pdcontact 62 -517 62 -517 1 anda1n
rlabel polycontact 96 -532 96 -532 1 anda1n
rlabel pdcontact 106 -517 106 -517 1 outanda1
rlabel ndcontact 106 -559 106 -559 1 outanda1
rlabel polycontact 139 -581 139 -581 1 outanda1
rlabel pdcontact 62 -595 62 -595 1 anda2n
rlabel ndcontact 74 -634 74 -634 1 anda2n
rlabel ndiffusion 62 -634 62 -634 1 anda2m
rlabel polycontact 96 -612 96 -612 1 anda2n
rlabel pdcontact 106 -595 106 -595 1 outanda2
rlabel ndcontact 106 -637 106 -637 1 outanda2
rlabel polycontact 147 -588 147 -588 1 outanda2
rlabel pdcontact 62 -679 62 -679 1 andb1n
rlabel ndiffusion 62 -718 62 -718 1 andb1m
rlabel ndcontact 74 -718 74 -718 1 andb1n
rlabel polycontact 96 -694 96 -694 1 andb1n
rlabel pdcontact 106 -679 106 -679 1 outband1
rlabel ndcontact 106 -721 106 -721 1 outband1
rlabel polycontact 142 -743 142 -743 1 outband1
rlabel pdcontact 62 -757 62 -757 1 andb2n
rlabel polycontact 96 -774 96 -774 1 andb2n
rlabel ndcontact 74 -796 74 -796 1 andb2n
rlabel ndiffusion 62 -796 62 -796 1 andb2m
rlabel pdcontact 106 -757 106 -757 1 outband2
rlabel ndcontact 106 -799 106 -799 1 outband2
rlabel polycontact 150 -750 150 -750 1 outband2
rlabel pdcontact 62 -841 62 -841 1 andc1n
rlabel polycontact 96 -856 96 -856 1 andc1n
rlabel ndcontact 74 -880 74 -880 1 andc1n
rlabel ndiffusion 62 -880 62 -880 1 andc1m
rlabel pdcontact 106 -841 106 -841 1 outcand1
rlabel ndcontact 106 -883 106 -883 1 outcand1
rlabel polycontact 139 -905 139 -905 1 outcand1
rlabel pdcontact 62 -919 62 -919 1 andc2n
rlabel ndcontact 74 -958 74 -958 1 andc2n
rlabel polycontact 96 -936 96 -936 1 andc2n
rlabel ndiffusion 62 -958 62 -958 1 andc2m
rlabel ndcontact 106 -961 106 -961 1 outcand2
rlabel pdcontact 106 -919 106 -919 1 outcand2
rlabel polycontact 147 -912 147 -912 1 outcand2
rlabel polycontact 584 -640 584 -640 1 g0
rlabel polycontact 538 -569 538 -569 1 g0
rlabel pdcontact 423 -564 423 -564 1 c3_bar
rlabel ndcontact 423 -616 423 -616 1 c3_bar
rlabel ndcontact 405 -616 405 -616 1 c3_bar
rlabel polycontact 445 -587 445 -587 1 c3_bar
rlabel ndcontact 546 -909 546 -909 1 c3_bar1
rlabel pdcontact 546 -884 546 -884 1 c3_bar1
rlabel polycontact 573 -885 573 -885 1 c3_bar1
rlabel polycontact 572 -720 572 -720 1 c2_bar1
rlabel ndcontact 545 -744 545 -744 1 c2_bar1
rlabel pdcontact 545 -719 545 -719 1 c2_bar1
rlabel ndcontact -88 -1137 -88 -1137 1 b3
rlabel metal1 -84 -1105 -84 -1105 1 b3
rlabel pdcontact -88 -1078 -88 -1078 1 b3
rlabel polycontact -95 -1105 -95 -1105 1 b3_bar
rlabel ndcontact -108 -1134 -108 -1134 1 b3_bar
rlabel pdcontact -108 -1078 -108 -1078 1 b3_bar
rlabel polycontact -129 -1105 -129 -1105 1 b3b
rlabel pdcontact -145 -1078 -145 -1078 1 b3b
rlabel ndcontact -145 -1134 -145 -1134 1 b3b
rlabel ndiffusion -120 -1134 -120 -1134 1 b3m3
rlabel ndiffusion -158 -1134 -158 -1134 1 b3m2
rlabel polycontact -154 -1120 -154 -1120 1 b3a
rlabel ndcontact -183 -1137 -183 -1137 1 b3a
rlabel pdcontact -183 -1084 -183 -1084 1 b3a
rlabel pdiffusion -195 -1084 -195 -1084 1 b3m1
rlabel polycontact -204 -1105 -204 -1105 1 b3in
rlabel ndcontact -88 -1030 -88 -1030 1 a3
rlabel metal1 -84 -998 -84 -998 1 a3
rlabel pdcontact -88 -971 -88 -971 1 a3
rlabel ndcontact -108 -1027 -108 -1027 1 a3_bar
rlabel polycontact -95 -998 -95 -998 1 a3_bar
rlabel pdcontact -108 -971 -108 -971 1 a3_bar
rlabel polycontact -129 -998 -129 -998 1 a3b
rlabel ndcontact -145 -1027 -145 -1027 1 a3b
rlabel pdcontact -145 -971 -145 -971 1 a3b
rlabel polycontact -154 -1013 -154 -1013 1 a3a
rlabel ndcontact -183 -1030 -183 -1030 1 a3a
rlabel pdcontact -183 -977 -183 -977 1 a3a
rlabel polycontact -204 -998 -204 -998 1 a3in
rlabel ndiffusion -120 -1027 -120 -1027 1 a3m3
rlabel ndiffusion -158 -1027 -158 -1027 1 a3m2
rlabel pdiffusion -195 -977 -195 -977 1 a3m1
rlabel pdcontact -88 -864 -88 -864 1 b2
rlabel ndcontact -88 -923 -88 -923 1 b2
rlabel metal1 -84 -891 -84 -891 1 b2
rlabel polycontact -95 -891 -95 -891 1 b2_bar
rlabel pdcontact -108 -864 -108 -864 1 b2_bar
rlabel ndcontact -108 -920 -108 -920 1 b2_bar
rlabel ndiffusion -120 -920 -120 -920 1 b2m3
rlabel polycontact -129 -891 -129 -891 1 b2b
rlabel ndcontact -145 -920 -145 -920 1 b2b
rlabel pdcontact -145 -864 -145 -864 1 b2b
rlabel polycontact -154 -906 -154 -906 1 b2a
rlabel ndcontact -183 -923 -183 -923 1 b2a
rlabel pdcontact -183 -870 -183 -870 1 b2a
rlabel polycontact -204 -891 -204 -891 1 b2in
rlabel ndiffusion -158 -920 -158 -920 1 b2m2
rlabel pdiffusion -195 -870 -195 -870 1 b2m1
rlabel pdcontact -88 -757 -88 -757 1 a2
rlabel ndcontact -88 -816 -88 -816 1 a2
rlabel metal1 -84 -784 -84 -784 1 a2
rlabel pdcontact -108 -757 -108 -757 1 a2_bar
rlabel ndcontact -108 -813 -108 -813 1 a2_bar
rlabel polycontact -95 -784 -95 -784 1 a2_bar
rlabel polycontact -129 -784 -129 -784 1 a2b
rlabel pdcontact -145 -757 -145 -757 1 a2b
rlabel ndcontact -145 -813 -145 -813 1 a2b
rlabel polycontact -154 -799 -154 -799 1 a2a
rlabel pdcontact -183 -763 -183 -763 1 a2a
rlabel ndcontact -183 -816 -183 -816 1 a2a
rlabel polycontact -204 -784 -204 -784 1 a2in
rlabel ndiffusion -120 -813 -120 -813 1 a2m3
rlabel ndiffusion -158 -813 -158 -813 1 a2m2
rlabel pdiffusion -195 -763 -195 -763 1 a2m1
rlabel pdcontact -88 -650 -88 -650 1 b1
rlabel ndcontact -88 -709 -88 -709 1 b1
rlabel metal1 -84 -677 -84 -677 1 b1
rlabel polycontact -95 -677 -95 -677 1 b1_bar
rlabel pdcontact -108 -650 -108 -650 1 b1_bar
rlabel ndcontact -108 -706 -108 -706 1 b1_bar
rlabel polycontact -129 -677 -129 -677 1 b1b
rlabel pdcontact -145 -650 -145 -650 1 b1b
rlabel ndcontact -145 -706 -145 -706 1 b1b
rlabel ndcontact -183 -709 -183 -709 1 b1a
rlabel polycontact -154 -692 -154 -692 1 b1a
rlabel pdcontact -183 -656 -183 -656 1 b1a
rlabel ndiffusion -120 -706 -120 -706 1 b1m3
rlabel ndiffusion -158 -706 -158 -706 1 b1m2
rlabel pdiffusion -195 -656 -195 -656 1 b1m1
rlabel pdcontact -88 -543 -88 -543 1 a1
rlabel metal1 -84 -570 -84 -570 1 a1
rlabel ndcontact -88 -602 -88 -602 1 a1
rlabel polycontact -95 -570 -95 -570 1 a1_bar
rlabel pdcontact -108 -543 -108 -543 1 a1_bar
rlabel ndcontact -108 -599 -108 -599 1 a1_bar
rlabel polycontact -129 -570 -129 -570 1 a1b
rlabel ndcontact -145 -599 -145 -599 1 a1b
rlabel pdcontact -145 -543 -145 -543 1 a1b
rlabel polycontact -154 -585 -154 -585 1 a1a
rlabel pdcontact -183 -549 -183 -549 1 a1a
rlabel ndcontact -183 -602 -183 -602 1 a1a
rlabel polycontact -204 -570 -204 -570 1 a1in
rlabel ndiffusion -120 -599 -120 -599 1 a1m3
rlabel ndiffusion -157 -599 -157 -599 1 a1m2
rlabel pdiffusion -195 -549 -195 -549 1 a1m1
rlabel ndcontact -88 -495 -88 -495 1 b0
rlabel pdcontact -88 -436 -88 -436 1 b0
rlabel metal1 -84 -463 -84 -463 1 b0
rlabel pdcontact -108 -436 -108 -436 1 b0_bar
rlabel polycontact -95 -463 -95 -463 1 b0_bar
rlabel ndcontact -108 -492 -108 -492 1 b0_bar
rlabel ndiffusion -120 -492 -120 -492 1 b0m3
rlabel pdcontact -145 -436 -145 -436 1 b0b
rlabel polycontact -129 -463 -129 -463 1 b0b
rlabel ndcontact -145 -492 -145 -492 1 b0b
rlabel ndiffusion -158 -492 -158 -492 1 b0m2
rlabel polycontact -154 -478 -154 -478 1 b0a
rlabel ndcontact -183 -495 -183 -495 1 b0a
rlabel pdcontact -183 -442 -183 -442 1 b0a
rlabel pdiffusion -195 -442 -195 -442 1 b0m1
rlabel polycontact -204 -463 -204 -463 1 b0in
rlabel pdcontact -88 -329 -88 -329 1 a0
rlabel metal1 -84 -356 -84 -356 1 a0
rlabel pdcontact -108 -329 -108 -329 1 a0_bar
rlabel polycontact -95 -356 -95 -356 1 a0_bar
rlabel ndcontact -88 -388 -88 -388 1 a0
rlabel ndcontact -108 -385 -108 -385 1 a0_bar
rlabel polycontact -129 -356 -129 -356 1 a0b
rlabel ndiffusion -120 -385 -120 -385 1 a0m3
rlabel pdcontact -145 -329 -145 -329 1 a0b
rlabel ndcontact -145 -385 -145 -385 1 a0b
rlabel ndiffusion -158 -385 -158 -385 1 a0m2
rlabel polycontact -154 -371 -154 -371 1 a0a
rlabel ndcontact -183 -388 -183 -388 1 a0a
rlabel pdcontact -183 -335 -183 -335 1 a0a
rlabel polycontact -204 -356 -204 -356 1 a0in
rlabel pdiffusion -195 -335 -195 -335 1 a0m1
rlabel ndcontact -108 -278 -108 -278 1 c0_bar
rlabel pdcontact -108 -222 -108 -222 1 c0_bar
rlabel polycontact -95 -249 -95 -249 1 c0_bar
rlabel ndcontact -88 -281 -88 -281 1 c0
rlabel metal1 -84 -249 -84 -249 1 c0
rlabel pdcontact -88 -222 -88 -222 1 c0
rlabel ndiffusion -120 -278 -120 -278 1 cinm3
rlabel polycontact -129 -249 -129 -249 1 cinb
rlabel ndcontact -145 -278 -145 -278 1 cinb
rlabel pdcontact -145 -222 -145 -222 1 cinb
rlabel ndiffusion -158 -278 -158 -278 1 cinm2
rlabel polycontact -154 -264 -154 -264 1 cino1
rlabel ndcontact -183 -281 -183 -281 1 cino1
rlabel pdcontact -183 -228 -183 -228 1 cino1
rlabel pdiffusion -195 -228 -195 -228 1 cinm
rlabel polycontact -204 -249 -204 -249 1 cin
rlabel polycontact -166 -249 -166 -249 1 CLK
rlabel polycontact -117 -256 -117 -256 1 CLK
rlabel polycontact -192 -256 -192 -256 1 CLK
rlabel pdcontact -96 -222 -96 -222 1 vdd
rlabel ndcontact -96 -281 -96 -281 1 gnd
rlabel pdcontact -132 -222 -132 -222 1 vdd
rlabel ndcontact -132 -278 -132 -278 1 gnd
rlabel pdcontact -169 -222 -169 -222 1 vdd
rlabel ndcontact -169 -278 -169 -278 1 gnd
rlabel pdcontact -207 -228 -207 -228 1 vdd
rlabel metal1 -139 -290 -139 -290 1 gnd
rlabel ndcontact -207 -281 -207 -281 1 gnd
rlabel metal1 -154 -209 -154 -209 5 VDD
rlabel polycontact -166 -356 -166 -356 1 CLK
rlabel polycontact -117 -363 -117 -363 1 CLK
rlabel polycontact -192 -363 -192 -363 1 CLK
rlabel pdcontact -96 -329 -96 -329 1 vdd
rlabel ndcontact -96 -388 -96 -388 1 gnd
rlabel pdcontact -132 -329 -132 -329 1 vdd
rlabel ndcontact -132 -385 -132 -385 1 gnd
rlabel pdcontact -169 -329 -169 -329 1 vdd
rlabel ndcontact -169 -385 -169 -385 1 gnd
rlabel pdcontact -207 -335 -207 -335 1 vdd
rlabel metal1 -139 -397 -139 -397 1 gnd
rlabel ndcontact -207 -388 -207 -388 1 gnd
rlabel metal1 -154 -316 -154 -316 5 VDD
rlabel polycontact -166 -463 -166 -463 1 CLK
rlabel polycontact -117 -470 -117 -470 1 CLK
rlabel polycontact -192 -470 -192 -470 1 CLK
rlabel pdcontact -96 -436 -96 -436 1 vdd
rlabel ndcontact -96 -495 -96 -495 1 gnd
rlabel pdcontact -132 -436 -132 -436 1 vdd
rlabel ndcontact -132 -492 -132 -492 1 gnd
rlabel pdcontact -169 -436 -169 -436 1 vdd
rlabel ndcontact -169 -492 -169 -492 1 gnd
rlabel pdcontact -207 -442 -207 -442 1 vdd
rlabel metal1 -139 -504 -139 -504 1 gnd
rlabel ndcontact -207 -495 -207 -495 1 gnd
rlabel metal1 -154 -423 -154 -423 5 VDD
rlabel polycontact -166 -570 -166 -570 1 CLK
rlabel polycontact -117 -577 -117 -577 1 CLK
rlabel polycontact -192 -577 -192 -577 1 CLK
rlabel pdcontact -96 -543 -96 -543 1 vdd
rlabel ndcontact -96 -602 -96 -602 1 gnd
rlabel pdcontact -132 -543 -132 -543 1 vdd
rlabel ndcontact -132 -599 -132 -599 1 gnd
rlabel pdcontact -169 -543 -169 -543 1 vdd
rlabel ndcontact -169 -599 -169 -599 1 gnd
rlabel pdcontact -207 -549 -207 -549 1 vdd
rlabel metal1 -139 -611 -139 -611 1 gnd
rlabel ndcontact -207 -602 -207 -602 1 gnd
rlabel metal1 -154 -530 -154 -530 5 VDD
rlabel polycontact -166 -677 -166 -677 1 CLK
rlabel polycontact -117 -684 -117 -684 1 CLK
rlabel polycontact -192 -684 -192 -684 1 CLK
rlabel pdcontact -96 -650 -96 -650 1 vdd
rlabel ndcontact -96 -709 -96 -709 1 gnd
rlabel pdcontact -132 -650 -132 -650 1 vdd
rlabel ndcontact -132 -706 -132 -706 1 gnd
rlabel pdcontact -169 -650 -169 -650 1 vdd
rlabel ndcontact -169 -706 -169 -706 1 gnd
rlabel pdcontact -207 -656 -207 -656 1 vdd
rlabel metal1 -139 -718 -139 -718 1 gnd
rlabel ndcontact -207 -709 -207 -709 1 gnd
rlabel metal1 -154 -637 -154 -637 5 VDD
rlabel polycontact -166 -784 -166 -784 1 CLK
rlabel polycontact -117 -791 -117 -791 1 CLK
rlabel polycontact -192 -791 -192 -791 1 CLK
rlabel pdcontact -96 -757 -96 -757 1 vdd
rlabel ndcontact -96 -816 -96 -816 1 gnd
rlabel pdcontact -132 -757 -132 -757 1 vdd
rlabel ndcontact -132 -813 -132 -813 1 gnd
rlabel pdcontact -169 -757 -169 -757 1 vdd
rlabel ndcontact -169 -813 -169 -813 1 gnd
rlabel pdcontact -207 -763 -207 -763 1 vdd
rlabel metal1 -139 -825 -139 -825 1 gnd
rlabel ndcontact -207 -816 -207 -816 1 gnd
rlabel metal1 -154 -744 -154 -744 5 VDD
rlabel polycontact -166 -891 -166 -891 1 CLK
rlabel polycontact -117 -898 -117 -898 1 CLK
rlabel polycontact -192 -898 -192 -898 1 CLK
rlabel pdcontact -96 -864 -96 -864 1 vdd
rlabel ndcontact -96 -923 -96 -923 1 gnd
rlabel pdcontact -132 -864 -132 -864 1 vdd
rlabel ndcontact -132 -920 -132 -920 1 gnd
rlabel pdcontact -169 -864 -169 -864 1 vdd
rlabel ndcontact -169 -920 -169 -920 1 gnd
rlabel pdcontact -207 -870 -207 -870 1 vdd
rlabel metal1 -139 -932 -139 -932 1 gnd
rlabel ndcontact -207 -923 -207 -923 1 gnd
rlabel metal1 -154 -851 -154 -851 5 VDD
rlabel polycontact -166 -998 -166 -998 1 CLK
rlabel polycontact -117 -1005 -117 -1005 1 CLK
rlabel polycontact -192 -1005 -192 -1005 1 CLK
rlabel pdcontact -96 -971 -96 -971 1 vdd
rlabel ndcontact -96 -1030 -96 -1030 1 gnd
rlabel pdcontact -132 -971 -132 -971 1 vdd
rlabel ndcontact -132 -1027 -132 -1027 1 gnd
rlabel pdcontact -169 -971 -169 -971 1 vdd
rlabel ndcontact -169 -1027 -169 -1027 1 gnd
rlabel pdcontact -207 -977 -207 -977 1 vdd
rlabel metal1 -139 -1039 -139 -1039 1 gnd
rlabel ndcontact -207 -1030 -207 -1030 1 gnd
rlabel metal1 -154 -958 -154 -958 5 VDD
rlabel polycontact -166 -1105 -166 -1105 1 CLK
rlabel polycontact -117 -1112 -117 -1112 1 CLK
rlabel polycontact -192 -1112 -192 -1112 1 CLK
rlabel pdcontact -96 -1078 -96 -1078 1 vdd
rlabel ndcontact -96 -1137 -96 -1137 1 gnd
rlabel pdcontact -132 -1078 -132 -1078 1 vdd
rlabel ndcontact -132 -1134 -132 -1134 1 gnd
rlabel pdcontact -169 -1078 -169 -1078 1 vdd
rlabel ndcontact -169 -1134 -169 -1134 1 gnd
rlabel pdcontact -207 -1084 -207 -1084 1 vdd
rlabel metal1 -139 -1146 -139 -1146 1 gnd
rlabel ndcontact -207 -1137 -207 -1137 1 gnd
rlabel metal1 -154 -1065 -154 -1065 5 VDD
rlabel ndcontact 907 -940 907 -940 1 s3f
rlabel metal1 911 -908 911 -908 7 s3f
rlabel pdcontact 907 -881 907 -881 1 s3f
rlabel ndiffusion 875 -937 875 -937 1 s3m3
rlabel polycontact 866 -908 866 -908 1 s3b
rlabel pdcontact 850 -881 850 -881 1 s3b
rlabel ndcontact 850 -937 850 -937 1 s3b
rlabel ndiffusion 838 -937 838 -937 1 s3m2
rlabel polycontact 841 -923 841 -923 1 s3a
rlabel ndcontact 812 -940 812 -940 1 s3a
rlabel pdcontact 812 -887 812 -887 1 s3a
rlabel pdiffusion 800 -887 800 -887 1 s3m1
rlabel polycontact 791 -908 791 -908 1 s3
rlabel metal1 841 -654 841 -654 5 VDD
rlabel ndcontact 788 -726 788 -726 1 gnd
rlabel metal1 856 -735 856 -735 1 gnd
rlabel pdcontact 788 -673 788 -673 1 vdd
rlabel ndcontact 826 -723 826 -723 1 gnd
rlabel pdcontact 826 -667 826 -667 1 vdd
rlabel ndcontact 863 -723 863 -723 1 gnd
rlabel pdcontact 863 -667 863 -667 1 vdd
rlabel ndcontact 899 -726 899 -726 1 gnd
rlabel pdcontact 899 -667 899 -667 1 vdd
rlabel polycontact 803 -701 803 -701 1 CLK
rlabel polycontact 878 -701 878 -701 1 CLK
rlabel polycontact 829 -694 829 -694 1 CLK
rlabel pdcontact 907 -774 907 -774 1 s2f
rlabel metal1 911 -801 911 -801 7 s2f
rlabel ndcontact 907 -833 907 -833 1 s2f
rlabel ndiffusion 875 -830 875 -830 1 s2m3
rlabel polycontact 866 -801 866 -801 1 s2b
rlabel ndcontact 850 -830 850 -830 1 s2b
rlabel pdcontact 850 -774 850 -774 1 s2b
rlabel ndiffusion 837 -830 837 -830 1 s2m2
rlabel polycontact 841 -816 841 -816 1 s2a
rlabel ndcontact 812 -833 812 -833 1 s2a
rlabel pdcontact 812 -780 812 -780 1 s2a
rlabel pdiffusion 800 -780 800 -780 1 s2m1
rlabel polycontact 791 -801 791 -801 1 s2
rlabel polycontact 829 -801 829 -801 1 CLK
rlabel polycontact 878 -808 878 -808 1 CLK
rlabel polycontact 803 -808 803 -808 1 CLK
rlabel pdcontact 899 -774 899 -774 1 vdd
rlabel ndcontact 899 -833 899 -833 1 gnd
rlabel pdcontact 863 -774 863 -774 1 vdd
rlabel ndcontact 863 -830 863 -830 1 gnd
rlabel pdcontact 826 -774 826 -774 1 vdd
rlabel ndcontact 826 -830 826 -830 1 gnd
rlabel pdcontact 788 -780 788 -780 1 vdd
rlabel metal1 856 -842 856 -842 1 gnd
rlabel ndcontact 788 -833 788 -833 1 gnd
rlabel metal1 841 -761 841 -761 5 VDD
rlabel pdcontact 907 -560 907 -560 1 s1f
rlabel ndcontact 907 -619 907 -619 1 s1f
rlabel metal1 911 -587 911 -587 7 s1f
rlabel ndiffusion 875 -616 875 -616 1 s1m3
rlabel polycontact 866 -587 866 -587 1 s1b
rlabel ndiffusion 837 -616 837 -616 1 s1m2
rlabel ndcontact 850 -616 850 -616 1 s1b
rlabel pdcontact 850 -560 850 -560 1 s1b
rlabel polycontact 841 -602 841 -602 1 s1a
rlabel ndcontact 812 -619 812 -619 1 s1a
rlabel pdcontact 812 -566 812 -566 1 s1a
rlabel polycontact 791 -587 791 -587 1 s1
rlabel pdiffusion 800 -566 800 -566 1 s1m1
rlabel ndcontact 907 -512 907 -512 1 s0f
rlabel pdcontact 907 -453 907 -453 1 s0f
rlabel metal1 911 -480 911 -480 7 s0f
rlabel ndiffusion 875 -509 875 -509 1 s0m3
rlabel polycontact 866 -480 866 -480 1 s0b
rlabel pdcontact 850 -453 850 -453 1 s0b
rlabel ndcontact 850 -509 850 -509 1 s0b
rlabel ndiffusion 837 -509 837 -509 1 s0m2
rlabel polycontact 841 -495 841 -495 1 s0a
rlabel ndcontact 812 -512 812 -512 1 s0a
rlabel pdcontact 812 -459 812 -459 1 s0a
rlabel pdiffusion 800 -459 800 -459 1 s0m1
rlabel polycontact 791 -480 791 -480 1 s0
rlabel polycontact 829 -480 829 -480 1 CLK
rlabel polycontact 878 -487 878 -487 1 CLK
rlabel polycontact 803 -487 803 -487 1 CLK
rlabel pdcontact 899 -453 899 -453 1 vdd
rlabel ndcontact 899 -512 899 -512 1 gnd
rlabel pdcontact 863 -453 863 -453 1 vdd
rlabel ndcontact 863 -509 863 -509 1 gnd
rlabel pdcontact 826 -453 826 -453 1 vdd
rlabel ndcontact 826 -509 826 -509 1 gnd
rlabel pdcontact 788 -459 788 -459 1 vdd
rlabel metal1 856 -521 856 -521 1 gnd
rlabel ndcontact 788 -512 788 -512 1 gnd
rlabel metal1 841 -440 841 -440 5 VDD
rlabel polycontact 829 -587 829 -587 1 CLK
rlabel polycontact 878 -594 878 -594 1 CLK
rlabel polycontact 803 -594 803 -594 1 CLK
rlabel pdcontact 899 -560 899 -560 1 vdd
rlabel ndcontact 899 -619 899 -619 1 gnd
rlabel pdcontact 863 -560 863 -560 1 vdd
rlabel ndcontact 863 -616 863 -616 1 gnd
rlabel pdcontact 826 -560 826 -560 1 vdd
rlabel ndcontact 826 -616 826 -616 1 gnd
rlabel pdcontact 788 -566 788 -566 1 vdd
rlabel metal1 856 -628 856 -628 1 gnd
rlabel ndcontact 788 -619 788 -619 1 gnd
rlabel metal1 841 -547 841 -547 5 VDD
rlabel polycontact 829 -908 829 -908 1 CLK
rlabel polycontact 878 -915 878 -915 1 CLK
rlabel polycontact 803 -915 803 -915 1 CLK
rlabel pdcontact 899 -881 899 -881 1 vdd
rlabel ndcontact 899 -940 899 -940 1 gnd
rlabel pdcontact 863 -881 863 -881 1 vdd
rlabel ndcontact 863 -937 863 -937 1 gnd
rlabel pdcontact 826 -881 826 -881 1 vdd
rlabel ndcontact 826 -937 826 -937 1 gnd
rlabel pdcontact 788 -887 788 -887 1 vdd
rlabel metal1 856 -949 856 -949 1 gnd
rlabel ndcontact 788 -940 788 -940 1 gnd
rlabel metal1 841 -868 841 -868 5 VDD
rlabel polycontact 791 -694 791 -694 1 cout
rlabel pdiffusion 800 -673 800 -673 1 coutm1
rlabel pdcontact 812 -673 812 -673 1 couta
rlabel ndcontact 812 -726 812 -726 1 couta
rlabel polycontact 841 -709 841 -709 1 couta
rlabel ndiffusion 838 -723 838 -723 1 coutm2
rlabel ndcontact 850 -723 850 -723 1 coutb
rlabel pdcontact 850 -667 850 -667 1 coutb
rlabel polycontact 866 -694 866 -694 1 coutb
rlabel ndiffusion 875 -723 875 -723 1 coutm3
rlabel metal1 911 -694 911 -694 1 coutf
rlabel pdcontact 907 -667 907 -667 1 coutf
rlabel ndcontact 907 -726 907 -726 1 coutf
rlabel polycontact -204 -677 -204 -677 1 b1in
rlabel polycontact 900 -694 900 -694 1 coutf_bar
rlabel pdcontact 887 -667 887 -667 1 coutf_bar
rlabel ndcontact 887 -723 887 -723 1 coutf_bar
rlabel pdcontact 887 -881 887 -881 1 s3f_bar
rlabel polycontact 900 -908 900 -908 1 s3f_bar
rlabel ndcontact 887 -937 887 -937 1 s3f_bar
rlabel ndcontact 887 -830 887 -830 1 s2f_bar
rlabel polycontact 900 -801 900 -801 1 s2f_bar
rlabel pdcontact 887 -774 887 -774 1 s2f_bar
rlabel ndcontact 887 -616 887 -616 1 s1f_bar
rlabel polycontact 900 -587 900 -587 1 s1f_bar
rlabel pdcontact 887 -560 887 -560 1 s1f_bar
rlabel ndcontact 887 -509 887 -509 1 s0f_bar
rlabel polycontact 900 -480 900 -480 1 s0f_bar
rlabel pdcontact 887 -453 887 -453 1 s0f_bar
<< end >>
